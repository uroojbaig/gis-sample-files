WKT,nameenglis,namearabic
"POLYGON ((58.0431701843931 23.4338248491112,57.9829898357381 23.4511725532561,57.9329829022871 23.4386300436554,57.925316766388 23.3997308309108,57.9295815083327 23.3806596380139,57.9243487084833 23.3694872861304,57.916959092147 23.3642090722159,57.915837256192 23.3553928613188,57.9066179016667 23.3483742717905,57.8898206922342 23.3300546725704,57.8809481580737 23.3291945398898,57.8609023186332 23.3114500597008,57.8568826250543 23.2990779171294,57.8730298085447 23.2887655491321,57.8631138000184 23.2548592225636,57.8239001949959 23.2337124500643,57.8212602440321 23.2106882094093,57.7911204071601 23.1456492286495,57.7873093976885 23.1426732898508,57.8066596186993 23.0904063239876,57.8083022097044 23.0859676153464,57.8299455517225 23.0838086593863,57.8391457747787 23.0702391263559,57.8618524629866 23.0715907244607,57.8712107864775 23.0638840694945,57.9154925011361 22.9906149628175,57.9487417858763 22.9915292475961,58.0003491763969 22.9826034811251,58.0177028761649 22.9763317560151,58.0227409928552 22.9672022340991,58.0371092498964 22.9757761136119,58.0381539627468 22.9961158970964,58.050671212359 23.003650618758,58.0835374477787 23.0189762118738,58.1254829253822 23.0172170316306,58.133590906604 23.0152727830984,58.1565137868418 23.0270438975178,58.1532019979003 23.0317526076623,58.1731934867358 23.03690684182,58.1698539614228 23.0463262691127,58.1915319942986 23.0557095492645,58.2012648035899 23.057314017844,58.2071401741386 23.0452263527211,58.2164037241019 23.052017045401,58.2303411890025 23.0523692863411,58.2346219933729 23.0642630120859,58.2564145969243 23.0755949816373,58.2952992662861 23.1191718154691,58.2711291315975 23.1723047973153,58.2617015721919 23.2191237709741,58.2209137728906 23.2313950833118,58.1899157345405 23.2791089074749,58.2129665615083 23.3210629188753,58.2132660634493 23.3426308256966,58.2068285201202 23.3500324030617,58.1676475320334 23.3374564703384,58.1544214135403 23.3369209299095,58.1305474514014 23.3687317329282,58.1263357888263 23.3766047862114,58.1123327711566 23.3733224629356,58.107161552849 23.3785767524944,58.1004858123198 23.364324459516,58.0773081063557 23.3606179020888,58.0740104403202 23.3891355451027,58.0431701843931 23.4338248491112))",Wilayat Samail,ولاية سمائل
"POLYGON ((57.6455202257619 23.5354355570249,57.6171772165899 23.551371610473,57.5973749106257 23.6152730935861,57.5330678986042 23.6091402681495,57.439983535349 23.5984343054152,57.4250709411323 23.6846540917876,57.3011150582473 23.6792457424469,57.2520651874765 23.6622722336727,57.1864983434453 23.61266944492,57.0909877707499 23.5647534226562,57.0360308316768 23.547668422976,57.0939741276902 23.5072933756842,57.0781111618808 23.4896179497523,57.0205122736929 23.4668760729069,57.0073974767621 23.4514719633033,57.0226635116953 23.4407785693073,57.0570409947282 23.4119548306984,57.0887326857516 23.3712242339003,57.0714485620544 23.3323487359329,57.0833631221438 23.3187908089929,57.1188660853235 23.3117556827149,57.1398326019131 23.3008695446255,57.1431457064386 23.2892888655115,57.1697322393798 23.27854889679,57.1853064160472 23.2620551664518,57.2023192742883 23.2620341670123,57.2642264609135 23.2448099945195,57.2707213717463 23.2326778043762,57.3285374807796 23.1957292645379,57.3698370217555 23.1793275261584,57.3948387209004 23.1814347312064,57.4322840535718 23.1643985881113,57.4429423167376 23.1553541340959,57.4632023306488 23.1509576653776,57.4746143952956 23.2364634735567,57.4915171624744 23.3111206638393,57.4967049496283 23.3244617048432,57.4876946539255 23.328408613135,57.4853412093886 23.3362842688902,57.4912445403521 23.3470107948915,57.503722876702 23.3491807255382,57.5709514673721 23.3872122866997,57.5726956960574 23.4100635263732,57.6196304705444 23.4279989122164,57.6231677438138 23.4852245904406,57.6455202257619 23.5354355570249))",Wilayat Ar Rustaq,ولاية الرستاق
"POLYGON ((57.5161348990359 23.8271157816073,57.4776408587699 23.8411150230172,57.4524703563945 23.8475820167646,57.4099710431765 23.860391799436,57.3664936889812 23.8712131665973,57.3362385595734 23.882056725215,57.3001806893868 23.8909473357666,57.2298030373389 23.9152306338502,57.1827794971621 23.9348198119062,57.1578851129231 23.9470759055079,57.1474968880666 23.9355898620164,57.1296629295869 23.8976201136269,57.1201831909695 23.8881978461004,57.1188784905335 23.8698430908918,57.129809038168 23.8544390712902,57.1606781928452 23.8274683318758,57.1631038455383 23.8209689799977,57.1609345582231 23.8092907268387,57.139077669174 23.7813307715453,57.1316368904858 23.7603178491982,57.1030783076364 23.6987133594241,57.0753594287983 23.6607331869273,57.0454157095675 23.655791147101,57.0416869804616 23.6308093871864,57.0909877707499 23.5647534226562,57.1864983434453 23.61266944492,57.2520651874765 23.6622722336727,57.3011150582473 23.6792457424469,57.4250709411323 23.6846540917876,57.4276118748351 23.7220477054225,57.4714990474708 23.7407654872652,57.4849876224037 23.7484042878331,57.5024876282156 23.7524071525977,57.5144974943696 23.7759008223496,57.5257107372459 23.782162136863,57.5386639773258 23.8030843883924,57.5181268104177 23.812849128255,57.5161348990359 23.8271157816073))",Wilayat As Suwayq,ولاية السويق
"POLYGON ((58.4785878338926 23.5598591517219,58.4766925809497 23.5734491991809,58.4912989118572 23.5791503096642,58.4898878192365 23.589275956937,58.4929588753045 23.5999161967475,58.4927305258314 23.6116347800732,58.4728614934133 23.6133441829714,58.4670827744354 23.6193216581268,58.453002234089 23.6130725933114,58.4215704826534 23.6056869267545,58.3904837714574 23.6036595352615,58.3692957970843 23.6056234652235,58.3393223641763 23.6057442119843,58.3283968131764 23.607419917078,58.3328655109609 23.60384345311,58.3292600413018 23.5920485793623,58.3168617203465 23.5894247011142,58.3179138970369 23.5810202348409,58.3260043773073 23.581991935827,58.3252994210079 23.5726759867235,58.3095448188354 23.554993277225,58.3061376362758 23.5470225443403,58.3056666946116 23.5250557923381,58.2983300951141 23.505210001385,58.2888306864344 23.5070821369266,58.2827956265455 23.5159758443596,58.2766744789048 23.5160261574616,58.2704215541234 23.5023410168578,58.2697771875059 23.4839829037692,58.2450239112885 23.4543713335279,58.251585954932 23.4271185147935,58.2669696902108 23.4189257150644,58.2826059172647 23.4007841401843,58.3065872602882 23.3785487103259,58.3103629333383 23.3689490051002,58.33321616107 23.3725671854633,58.3388002677574 23.3780505805348,58.3403933529886 23.3888910418597,58.3652856508999 23.3836433427898,58.3680152368453 23.3961198668439,58.3621610726008 23.4038634221309,58.3724129657688 23.4058767426011,58.3837051251011 23.4222048250889,58.387283216214 23.4426466474039,58.3950576436073 23.4530376044491,58.3898726680574 23.4608157442214,58.3827508147272 23.4600481840032,58.3768679805197 23.4656498501201,58.3905911362266 23.4833654667954,58.4026491998197 23.4928844877897,58.4070052496607 23.5040030162455,58.4177931720052 23.5124823457155,58.4243949104989 23.5290841645231,58.4437528850059 23.5353718803566,58.4578004998565 23.54815045086,58.4785878338926 23.5598591517219))",Wilayat Bawshar,ولاية بوشر
"POLYGON ((58.0816830738052 23.5628765732803,58.0535001300214 23.5821584504815,58.0278021330441 23.5926053969556,58.0085388161426 23.5919040394889,57.9923532749528 23.5821922588092,57.968495634177 23.5347928616926,57.9361421317924 23.5058871782189,57.9016338482612 23.4924878393072,57.8660666755163 23.4527460693535,57.8586918902918 23.4385241690305,57.8302605652216 23.4323536724689,57.8243247798967 23.4149544982799,57.8180735031818 23.4183459874182,57.8058213908944 23.3895368130702,57.7932180207431 23.3860179162521,57.7804870542067 23.3878336634047,57.758721882507 23.3811127742887,57.7497334593949 23.3673590061664,57.7461373289791 23.3564111953012,57.7331126660347 23.3281278480357,57.7439987874604 23.2940925465078,57.772626351413 23.2823209555063,57.7663878817527 23.2615415882556,57.7750962252959 23.2476504281704,57.8048327352544 23.2320976161454,57.8049344421057 23.2281594113771,57.7787622281834 23.2200677526451,57.778896575811 23.2013043648511,57.7946759110232 23.1929258729439,57.7943290199731 23.1841919150161,57.7833472852815 23.1839392207117,57.7605033068958 23.1897274205329,57.7496274534921 23.181199460108,57.7545966577451 23.1638734728634,57.7474633055432 23.1574932986436,57.739834862516 23.1611584521895,57.7277678477971 23.1877827064313,57.7125591842319 23.1944733934047,57.7026939609394 23.2111053587901,57.6797891712134 23.2430082488565,57.6800066226663 23.2561449307578,57.6711841716663 23.3244024499799,57.693339536708 23.3292305007318,57.7238832118698 23.3459422534408,57.7284412401867 23.3521868562222,57.7404375923741 23.3938964461694,57.7403484338001 23.431360497841,57.7839072160613 23.4696439618809,57.7810608223676 23.4991788719302,57.7539008111138 23.5186070512728,57.708975943153 23.5397030777987,57.6965770727845 23.533797548686,57.6904054401984 23.5383397873566,57.6455202257619 23.5354355570249,57.6231677438138 23.4852245904406,57.6196304705444 23.4279989122164,57.6772612147052 23.406356455679,57.6710080449743 23.3645947976413,57.6555570780715 23.3554425652139,57.6218100512967 23.3760957464374,57.6010671038242 23.3525896330669,57.587816384524 23.3518179041022,57.5872014824808 23.3469567426927,57.5982317373016 23.3429859883415,57.6024355784288 23.3316645223308,57.6304136740542 23.3311386374251,57.6311901993938 23.3048811889991,57.6273497346466 23.2813151526135,57.638398386187 23.2520699210896,57.6254265928873 23.2274356581371,57.6608193563938 23.1899296820924,57.6802499238108 23.1790999749658,57.6951789063901 23.1562320103669,57.7209750331172 23.1621620425334,57.7194516355502 23.1320575903342,57.7351207964276 23.1189604059127,57.7574451686242 23.1193450072182,57.7873093976885 23.1426732898508,57.7911204071601 23.1456492286495,57.8212602440321 23.2106882094093,57.8239001949959 23.2337124500643,57.8631138000184 23.2548592225636,57.8730298085447 23.2887655491321,57.8568826250543 23.2990779171294,57.8609023186332 23.3114500597008,57.8809481580737 23.3291945398898,57.8898206922342 23.3300546725704,57.9066179016667 23.3483742717905,57.915837256192 23.3553928613188,57.916959092147 23.3642090722159,57.9243487084833 23.3694872861304,57.9295815083327 23.3806596380139,57.925316766388 23.3997308309108,57.9329829022871 23.4386300436554,57.9829898357381 23.4511725532561,58.0431701843931 23.4338248491112,58.0609506795656 23.4743454336585,58.0609281457484 23.51297899983,58.0745994589962 23.5389658854337,58.0816830738052 23.5628765732803))",Wilayat Nakhal,ولاية نخل
"POLYGON ((58.3283968131764 23.607419917078,58.2901359282043 23.617953564596,58.2614054693189 23.6323613922161,58.2382816932107 23.6470598353386,58.2081411590203 23.6722751815208,58.1963069238491 23.6802592548253,58.1705721356672 23.6913342988481,58.1406834073912 23.701901960988,58.1148089248992 23.7091112441533,58.0931108395057 23.7132357836976,58.0687978254054 23.7135745793987,58.064149894467 23.7005440872851,58.0645524901368 23.6932460825867,58.0782011980285 23.690869463789,58.0778072695916 23.677126253309,58.0864536473341 23.6687285490993,58.0741977322513 23.6570822656575,58.0753441027865 23.6513799411948,58.0897699333467 23.6319932695804,58.0865196381516 23.6198687472315,58.0870370644335 23.6097311157798,58.0924556065835 23.6047573186043,58.0954386276463 23.5803891506245,58.0816830738052 23.5628765732803,58.0745994589962 23.5389658854337,58.0609281457484 23.51297899983,58.0766447333544 23.5007623240994,58.1497816159235 23.4946910270113,58.1632584525037 23.4784061494495,58.1835042052094 23.4733763968563,58.1881570766493 23.4748219797359,58.2303666073906 23.463611508124,58.2311261335369 23.4590350237451,58.2450239112885 23.4543713335279,58.2697771875059 23.4839829037692,58.2704215541234 23.5023410168578,58.2766744789048 23.5160261574616,58.2827956265455 23.5159758443596,58.2888306864344 23.5070821369266,58.2983300951141 23.505210001385,58.3056666946116 23.5250557923381,58.3061376362758 23.5470225443403,58.3095448188354 23.554993277225,58.3252994210079 23.5726759867235,58.3260043773073 23.581991935827,58.3179138970369 23.5810202348409,58.3168617203465 23.5894247011142,58.3292600413018 23.5920485793623,58.3328655109609 23.60384345311,58.3283968131764 23.607419917078))",Wilayat As Seeb,ولاية السيب
"POLYGON ((56.518024239392 23.8318598840931,56.4937435796985 23.8467042771889,56.4959760999532 23.8603478151807,56.4926251315816 23.8688848934993,56.4842043452951 23.8727917874405,56.4854548428578 23.8921986298928,56.4741337093871 23.9016581108768,56.4663178334335 23.9012920328476,56.4606808425383 23.9090062207439,56.4393659729854 23.9160925606266,56.4062985821457 23.9139597283266,56.3832749616439 23.9301834479269,56.4014576689634 23.9398592916329,56.3970739512362 23.9471403379448,56.3954714206649 23.9590334154566,56.3903805601555 23.9590132852871,56.3773207647941 23.9744963081262,56.366095289422 23.9764176849778,56.3450448348159 23.9724893199336,56.2952571303968 23.9737116853177,56.2954478619075 23.9359585150791,56.2864005821546 23.9275585527684,56.2726178035238 23.9251882218804,56.2692743201292 23.9064384579195,56.2589982613359 23.8942842976786,56.2367547401094 23.8921580531834,56.2134305195452 23.8615188307404,56.2158231775628 23.8395851025108,56.2297699399721 23.8308298589116,56.2342403376419 23.8330925220435,56.2421722466205 23.8230420799869,56.2488374706065 23.808087429152,56.2411652750836 23.7806692419272,56.2475284159249 23.7634072887298,56.2397553653449 23.7484125065191,56.2564615331136 23.7472341328859,56.2354568548735 23.7362054440295,56.2328727085248 23.7386767654326,56.2099418397722 23.7242124879435,56.1979556389328 23.6766060328896,56.2340465725023 23.6321142929766,56.3210002847985 23.6351132977603,56.3625740904484 23.6194679289197,56.4173878650064 23.5929912272189,56.4835728384993 23.5433607695525,56.5100036876417 23.5346996466029,56.5467828997703 23.5263592717704,56.556519705645 23.5312733936119,56.5829814820682 23.5354524437455,56.6041445054678 23.5582641288564,56.5868366595159 23.5756656117063,56.5769052839787 23.575272602902,56.5693422813295 23.5884351864717,56.5890205236688 23.6023614101895,56.5807482466519 23.6144081701142,56.599699150996 23.6236586706037,56.5927062729867 23.6474799627038,56.5659146553283 23.6589533195302,56.5669245366057 23.6774027928617,56.5900527862972 23.7167430648257,56.5673795941769 23.7551589952148,56.5498596450383 23.7831032543773,56.5411386378796 23.8173927328728,56.518024239392 23.8318598840931))",Wilayat Yanqul,ولاية ينقل
"POLYGON ((57.9923532749528 23.5821922588092,57.880732222366 23.5595300568129,57.8517497080017 23.5757797684817,57.7346941486798 23.5919576099111,57.7163510517146 23.5869053670187,57.6904054401984 23.5383397873566,57.6965770727845 23.533797548686,57.708975943153 23.5397030777987,57.7539008111138 23.5186070512728,57.7810608223676 23.4991788719302,57.7839072160613 23.4696439618809,57.7403484338001 23.431360497841,57.7404375923741 23.3938964461694,57.7284412401867 23.3521868562222,57.7238832118698 23.3459422534408,57.693339536708 23.3292305007318,57.6711841716663 23.3244024499799,57.6800066226663 23.2561449307578,57.6797891712134 23.2430082488565,57.7026939609394 23.2111053587901,57.7125591842319 23.1944733934047,57.7277678477971 23.1877827064313,57.739834862516 23.1611584521895,57.7474633055432 23.1574932986436,57.7545966577451 23.1638734728634,57.7496274534921 23.181199460108,57.7605033068958 23.1897274205329,57.7833472852815 23.1839392207117,57.7943290199731 23.1841919150161,57.7946759110232 23.1929258729439,57.778896575811 23.2013043648511,57.7787622281834 23.2200677526451,57.8049344421057 23.2281594113771,57.8048327352544 23.2320976161454,57.7750962252959 23.2476504281704,57.7663878817527 23.2615415882556,57.772626351413 23.2823209555063,57.7439987874604 23.2940925465078,57.7331126660347 23.3281278480357,57.7461373289791 23.3564111953012,57.7497334593949 23.3673590061664,57.758721882507 23.3811127742887,57.7804870542067 23.3878336634047,57.7932180207431 23.3860179162521,57.8058213908944 23.3895368130702,57.8180735031818 23.4183459874182,57.8243247798967 23.4149544982799,57.8302605652216 23.4323536724689,57.8586918902918 23.4385241690305,57.8660666755163 23.4527460693535,57.9016338482612 23.4924878393072,57.9361421317924 23.5058871782189,57.968495634177 23.5347928616926,57.9923532749528 23.5821922588092))",Wilayat Wadi Al Maawil,ولاية وادي المعاول
"POLYGON ((57.6290960608466 22.5949951799129,57.6233305381534 22.6412756038783,57.6453876407389 22.7071371972214,57.6862538015027 22.7665058858992,57.6957295848235 22.795006433185,57.6997756681934 22.8161933556045,57.7333744794623 22.8322430634833,57.732812946825 22.8845917339745,57.6963889938017 22.8772161150716,57.6572502949887 22.8731247677458,57.6291797833739 22.8571056698022,57.5999156353851 22.8302290877283,57.5648640386637 22.8283951376657,57.5554875179866 22.7780673765756,57.5290406914977 22.7482457803368,57.4789929840942 22.6862691275745,57.5110075378977 22.584367006355,57.5260935933885 22.5814276801781,57.5283106520874 22.5667773497906,57.5597431958942 22.5437727907137,57.6290960608466 22.5949951799129))",Wilayat Manah,ولاية منح
"POLYGON ((56.2952571303968 23.9737116853177,56.232149805596 23.9817689174369,56.1763086486729 24.0135549421218,56.0491477429145 24.0150770941752,56.0626717479292 23.9742479129458,56.0688203279901 23.9622188486238,56.0689328201332 23.9465518998928,56.0443963640888 23.9422538863052,55.9612248017993 23.8986878881513,56.0008001893264 23.8456139100185,56.0050295125467 23.8070601784067,56.001553811727 23.7843136991836,55.9916142425238 23.7192262102091,56.0981746644668 23.645972297091,56.0654059990687 23.6101384860241,56.053603006396 23.57587050602,56.0325694371101 23.5530913845379,56.0534724313316 23.5338590958004,56.0334187440128 23.4988186248187,56.0109662657225 23.4792860447887,56.1485011860388 23.4939850819043,56.1790339050576 23.4847705687005,56.2083120155417 23.4872800509741,56.2631127896109 23.4741173021943,56.4192742947264 23.3847977879979,56.4539275287672 23.3780416738995,56.4692526684279 23.3717531193742,56.4835895012901 23.3784306596902,56.5504869848093 23.355865940678,56.5576416640074 23.3636689257919,56.551349879102 23.3777749651719,56.5606982588578 23.3835663763382,56.5806829372253 23.3836212365197,56.5734298584468 23.4057963843117,56.5824543749168 23.4161975132628,56.5786542827293 23.4326171454959,56.5864089702656 23.4502206615106,56.5568653044212 23.4862639990812,56.5821823497219 23.5026692395139,56.5829814820682 23.5354524437455,56.556519705645 23.5312733936119,56.5467828997703 23.5263592717704,56.5100036876417 23.5346996466029,56.4835728384993 23.5433607695525,56.4173878650064 23.5929912272189,56.3625740904484 23.6194679289197,56.3210002847985 23.6351132977603,56.2340465725023 23.6321142929766,56.1979556389328 23.6766060328896,56.2099418397722 23.7242124879435,56.2328727085248 23.7386767654326,56.2354568548735 23.7362054440295,56.2564615331136 23.7472341328859,56.2397553653449 23.7484125065191,56.2475284159249 23.7634072887298,56.2411652750836 23.7806692419272,56.2488374706065 23.808087429152,56.2421722466205 23.8230420799869,56.2342403376419 23.8330925220435,56.2297699399721 23.8308298589116,56.2158231775628 23.8395851025108,56.2134305195452 23.8615188307404,56.2367547401094 23.8921580531834,56.2589982613359 23.8942842976786,56.2692743201292 23.9064384579195,56.2726178035238 23.9251882218804,56.2864005821546 23.9275585527684,56.2954478619075 23.9359585150791,56.2952571303968 23.9737116853177))",Wilayat Dank,ولاية ضنك
"POLYGON ((57.9487417858763 22.9915292475961,57.9154925011361 22.9906149628175,57.8712107864775 23.0638840694945,57.8618524629866 23.0715907244607,57.8391457747787 23.0702391263559,57.8299455517225 23.0838086593863,57.8083022097044 23.0859676153464,57.8066596186993 23.0904063239876,57.7368914189014 23.0069873825142,57.7131896224724 22.98712305299,57.6969033549002 22.9608448764559,57.7263447325872 22.9388771366702,57.7251716134998 22.9241789278708,57.732812946825 22.8845917339745,57.7333744794623 22.8322430634833,57.6997756681934 22.8161933556045,57.6957295848235 22.795006433185,57.6862538015027 22.7665058858992,57.6453876407389 22.7071371972214,57.6233305381534 22.6412756038783,57.6290960608466 22.5949951799129,57.6365977437997 22.5347363600622,57.6263304123396 22.4949944380171,57.632788068992 22.4868555899997,57.6306030942587 22.4726745201264,57.6377532544282 22.4596392336495,57.6512890758618 22.452293269284,57.6862719150105 22.4521483058827,57.7005195628586 22.4605613950939,57.7020623407205 22.4721822026744,57.6759015291704 22.4996876378843,57.6744523732107 22.5137949020557,57.90430268359 22.603321718951,57.9051693936022 22.6486938755621,57.9735638613173 22.7133353558484,57.981793276584 22.7329213130798,57.9924346854956 22.7889106780778,57.9559003499965 22.8165969614619,57.9771333974979 22.827669082908,57.98876770748 22.8318062014249,57.9948486747811 22.8428695972614,58.011027978084 22.8638078189266,57.9973263049985 22.8709042115709,57.994561339742 22.8844408048127,57.9869362174441 22.8967911833011,57.974654914508 22.9085171004933,57.9734289765502 22.9180215482237,57.9529666656578 22.9498597174323,57.9487417858763 22.9915292475961))",Wilayat Izki,ولاية إزكي
"POLYGON ((59.2331441681103 22.5035754938877,59.209772993222 22.4992422613091,59.1736786927296 22.4969741318787,59.161667340915 22.5001145713279,59.1389875293776 22.5111830453867,59.1222644869574 22.5226186661547,59.1141053700098 22.5251219985034,59.1083267021768 22.5355751168756,59.1025486189412 22.5393845043202,59.084405639777 22.542568859845,59.06591531823 22.5412204666424,59.0543471702845 22.5345872373995,59.0454142858277 22.5366605509862,59.0348121129839 22.5329279527467,59.0315736550743 22.5196971210314,59.0122723234739 22.5005336368078,58.9968437811539 22.4932466999841,58.9661038543778 22.4919330389927,58.9647240994262 22.4724170222006,58.9566149780496 22.4607669083376,58.9374234812086 22.4482378017567,58.9355697599668 22.4427522576202,58.9445792584638 22.4302514591467,58.964782559812 22.413483659937,58.9918883004013 22.3875105357664,59.0034754767876 22.3809426214505,59.0162964031917 22.3805023218107,59.0263228868264 22.3681118687284,59.0517012801913 22.3584025638822,59.0631964949916 22.3449178719158,59.0712199582506 22.3401651248328,59.0798828581025 22.328090374862,59.0887532777067 22.3229585335157,59.0837304493275 22.297115514141,59.0904368161967 22.2922986610043,59.1230013385636 22.2858527245142,59.1383302330333 22.2802186423179,59.1452985123342 22.2647310076705,59.1444649493334 22.2551908122804,59.1297383445964 22.2218177785633,59.1318951114234 22.2027054855092,59.1375507972597 22.195578730064,59.1600213253434 22.1862078935266,59.1669401856022 22.1698508772806,59.1856856200291 22.1696004975564,59.1969303456648 22.1755441300137,59.2106562390264 22.1760037594312,59.2158601768061 22.1720611443688,59.2310256614561 22.1496129056054,59.2389374010541 22.1541243755708,59.2451422807889 22.1509835288419,59.2580142259424 22.1350736069301,59.2704260923883 22.1446809004468,59.2808465370564 22.1787498499918,59.2894572809357 22.2004706007885,59.3015387876658 22.201413034494,59.3044401767764 22.2164279735702,59.3144777249982 22.2290339600684,59.3269375799301 22.2308584965844,59.3321725489509 22.2369168990017,59.3298661263579 22.2542333590579,59.3361026369146 22.2609335141734,59.3601192029617 22.2615139640533,59.3723040386607 22.2732994674986,59.3619937490122 22.2953287346222,59.3654952130732 22.3075770758188,59.3561132838648 22.318257011333,59.3433057583592 22.3265618482268,59.343344014509 22.3346578633936,59.331803076603 22.3477988559574,59.3182287640147 22.3557509258289,59.3180824112286 22.3651757600971,59.328521746056 22.3882097102626,59.3449064622558 22.3865278091828,59.3521537089643 22.3815539082376,59.363677211843 22.385906560427,59.3652619442479 22.3934340457156,59.3621676585898 22.4052806311723,59.3246002191719 22.421586697767,59.3038829206835 22.4403657172698,59.2915917184511 22.4568108319012,59.279635769476 22.4599665915565,59.2590362810292 22.4811541803344,59.2539131847511 22.4970177183618,59.2484920064373 22.4953034792113,59.2331441681103 22.5035754938877))",Wilayat Al Kamil Wa Al Wafi,ولاية الكامل والوافي
"POLYGON ((57.6951789063901 23.1562320103669,57.6802499238108 23.1790999749658,57.6608193563938 23.1899296820924,57.6254265928873 23.2274356581371,57.638398386187 23.2520699210896,57.6273497346466 23.2813151526135,57.6311901993938 23.3048811889991,57.6304136740542 23.3311386374251,57.6024355784288 23.3316645223308,57.5982317373016 23.3429859883415,57.5872014824808 23.3469567426927,57.587816384524 23.3518179041022,57.6010671038242 23.3525896330669,57.6218100512967 23.3760957464374,57.6555570780715 23.3554425652139,57.6710080449743 23.3645947976413,57.6772612147052 23.406356455679,57.6196304705444 23.4279989122164,57.5726956960574 23.4100635263732,57.5709514673721 23.3872122866997,57.503722876702 23.3491807255382,57.4912445403521 23.3470107948915,57.4853412093886 23.3362842688902,57.4876946539255 23.328408613135,57.4967049496283 23.3244617048432,57.4915171624744 23.3111206638393,57.4746143952956 23.2364634735567,57.4632023306488 23.1509576653776,57.4976552966017 23.164894661691,57.5043366156789 23.1817025339094,57.5411958732754 23.1793392438928,57.5932300375817 23.1679473606814,57.6053570126213 23.1545259142653,57.6148477758737 23.1610017117779,57.6254189111624 23.155427904989,57.6745225981536 23.1516538592947,57.6951789063901 23.1562320103669))",Wilayat Al Awabi,ولاية العوابي
"POLYGON ((58.5711442207629 23.6227946763361,58.563351552717 23.6367965638809,58.5408010225341 23.6318133571784,58.5345353177238 23.6336761850928,58.5176888988406 23.6310287113534,58.5097000618632 23.6345447383561,58.5029220355388 23.6452865311116,58.4917098840513 23.640480250819,58.480825421287 23.6316108405826,58.4794372338077 23.6251830356729,58.4670827744354 23.6193216581268,58.4728614934133 23.6133441829714,58.4927305258314 23.6116347800732,58.4929588753045 23.5999161967475,58.4898878192365 23.589275956937,58.4912989118572 23.5791503096642,58.4766925809497 23.5734491991809,58.4785878338926 23.5598591517219,58.4969936846236 23.5610351985743,58.500503170204 23.5521829012917,58.5136226772524 23.5516854953891,58.5170343842621 23.5663766990957,58.5252172268422 23.5713627841786,58.5367718596606 23.5636858498291,58.551664830817 23.5504210435053,58.5675521098307 23.5330811698927,58.5847219754276 23.5248036403525,58.5881597371589 23.5296156981414,58.5741984274628 23.5455022213126,58.575522086622 23.549053599282,58.592129813898 23.5416059320111,58.5900879017391 23.5507407849228,58.59321520152 23.5638480266928,58.5891973948299 23.5683230908684,58.5828037693415 23.5915039547983,58.5796017945865 23.592859512025,58.5778902394246 23.6133398207,58.5711442207629 23.6227946763361))",Wilayat Mutrah,ولاية مطرح
"POLYGON ((58.5847219754276 23.5248036403525,58.5675521098307 23.5330811698927,58.551664830817 23.5504210435053,58.5367718596606 23.5636858498291,58.5252172268422 23.5713627841786,58.5170343842621 23.5663766990957,58.5136226772524 23.5516854953891,58.500503170204 23.5521829012917,58.4969936846236 23.5610351985743,58.4785878338926 23.5598591517219,58.4578004998565 23.54815045086,58.4437528850059 23.5353718803566,58.4243949104989 23.5290841645231,58.4177931720052 23.5124823457155,58.4070052496607 23.5040030162455,58.4026491998197 23.4928844877897,58.3905911362266 23.4833654667954,58.3768679805197 23.4656498501201,58.3827508147272 23.4600481840032,58.3898726680574 23.4608157442214,58.3950576436073 23.4530376044491,58.387283216214 23.4426466474039,58.3837051251011 23.4222048250889,58.3724129657688 23.4058767426011,58.3621610726008 23.4038634221309,58.3680152368453 23.3961198668439,58.3652856508999 23.3836433427898,58.3403933529886 23.3888910418597,58.3388002677574 23.3780505805348,58.33321616107 23.3725671854633,58.3103629333383 23.3689490051002,58.3038883830302 23.3431774662158,58.3374742039902 23.3168859046639,58.3297494310354 23.3078768010933,58.340132360524 23.2711528432161,58.3609041939617 23.2660065714797,58.374533190659 23.2514838282314,58.3573732076725 23.2482179489343,58.3675820218537 23.2285720096729,58.38338684108 23.2164818301514,58.4064739240594 23.223063835773,58.4105742777666 23.2298573679404,58.4463689847575 23.2487806996584,58.455074654626 23.2154807835916,58.4897210743145 23.1912509287535,58.5110534888391 23.2078121959091,58.5662278435041 23.2181382244103,58.5760759733906 23.2066541371709,58.5719923704017 23.2022129480979,58.6130011825488 23.1617850176371,58.6252309641002 23.1557603258174,58.64993211387 23.1588424558009,58.6553744916942 23.1736400492165,58.6499532761094 23.181007638388,58.6411442251497 23.186115638809,58.6473923208393 23.1922022590651,58.6406000435988 23.2047749193978,58.641809496159 23.2158519148404,58.6376798841718 23.2244911371558,58.6442717592705 23.2304163790255,58.6529235647498 23.2294956102664,58.6570281828067 23.2362084829656,58.6551410075431 23.2577900360585,58.6515934640506 23.2599335263041,58.6486338107098 23.2767904015974,58.6510082979457 23.3072588722463,58.6568020714895 23.3267396812778,58.664326730758 23.3372300337437,58.638270257022 23.3436420579431,58.6414001474914 23.3630197984674,58.6344148283239 23.3710866482078,58.6206066818597 23.375935204278,58.6163729554265 23.384819937205,58.6243313918009 23.3902244983827,58.6172525205831 23.3967785347809,58.6255631213109 23.4028646495428,58.6226341876613 23.4118646205401,58.6345923660847 23.4214363764844,58.6495079369714 23.4293967135926,58.6541283952234 23.4377974934615,58.6568400938258 23.4552247486703,58.6538429551246 23.4770902163348,58.6608872950006 23.4817478351413,58.6621787776166 23.4975298828955,58.6472885230882 23.5030283020613,58.6337914657881 23.5046284533534,58.6284279137012 23.4991443029832,58.6207120472031 23.5016304521277,58.6066005917651 23.5112535927542,58.5973332833092 23.5218853266507,58.5847219754276 23.5248036403525))",Wilayat Al Amrat,ولاية العامرات
"POLYGON ((57.3372691882338 23.0484531624246,57.305522226557 23.042988511844,57.2814620539525 23.0499244595369,57.2886851535063 23.0763366620951,57.2891911653837 23.0878774519778,57.2755310663946 23.0880526681774,57.2723047629798 23.0967141213756,57.2531973483078 23.0924724660662,57.240914074945 23.0846407617468,57.227497793227 23.0793982517919,57.2258391415713 23.0592907027261,57.2068323656364 23.0519084230132,57.2043232994765 23.0456930534614,57.1866756932885 23.0365571568731,57.1594391046784 23.0322536277856,57.1500223538638 23.0281073518141,57.133868217636 23.0273300039486,57.1240471750004 23.0324255196848,57.1364830571854 23.0542347628224,57.15130461537 23.1103180353977,57.1385277083 23.1339107546882,57.1332066715746 23.1714850563445,57.1201727184826 23.1774571506577,57.115596605321 23.1883239420253,57.1054231819287 23.1900533313597,57.0966890710622 23.2007898116578,57.0779359578782 23.2145284396679,57.0244831848497 23.2001290237258,56.9590998319249 23.1836492792936,56.963560369944 23.1565015695223,56.9572868956513 23.1559383052667,56.9313781645423 23.16547803008,56.9299717622437 23.1456307864969,56.9574901031644 23.1163023606107,56.929415571604 23.0677135637285,56.9213929694591 23.062449641667,56.9130726674589 23.0488374384913,56.915082597034 23.0439311272938,56.931644107119 23.0400317235076,56.946484281847 23.0318274979794,56.9226550939765 22.962636479535,56.9348290737217 22.954366638528,56.9389730117577 22.9295652498818,56.9177720985311 22.9082105308374,56.9077768586653 22.8927282047229,56.8884489487416 22.8906727468172,56.8888055479081 22.8851274348799,56.8977012127194 22.8771171252853,56.8860982313042 22.859134377095,56.9053017778457 22.8303121139811,56.9392312277962 22.8031788424478,56.9525515667859 22.8082388722136,56.990301019235 22.7758529274121,56.9961539857765 22.7595632269188,56.9850586887522 22.7324124953675,56.9457195290254 22.7292208449242,56.8890389962391 22.7185187189212,56.8376363063073 22.6870180692113,56.7822537152524 22.6369585451552,56.7786437565569 22.6251572444698,56.7597455616434 22.5852141336849,56.7648775493956 22.5406902607666,56.7872951725845 22.5047701604025,56.7871135066467 22.487152246743,56.7977129778548 22.4806327363134,56.7986486023276 22.4717073038441,56.786940139017 22.4703368349447,56.7862432386579 22.4027187697778,56.7744479601071 22.3534560655595,56.7739113587372 22.3118855840309,56.762836778117 22.2940622063036,56.9182809820048 22.2559094318221,56.9515337082296 22.2472972381213,56.9842370853745 22.2412150931346,56.9986535579405 22.2411066630328,57.0038661237096 22.2665827974693,57.0045990750416 22.2921832595225,57.0174573355013 22.3061653155684,57.080678491111 22.3440863340711,57.1013375710192 22.4604857861491,57.1325869331343 22.4892925121657,57.1878978133028 22.4567076816885,57.2107083976502 22.4604932020885,57.2405508589168 22.4884784600897,57.3167473924131 22.5359146574757,57.3303610021942 22.5388399480485,57.3305893732544 22.543883273411,57.3420319232345 22.5505505785692,57.3648990594252 22.5558071468251,57.3800724845484 22.5631553882492,57.3875149441882 22.5594459308724,57.3832967815503 22.5502026199542,57.5130171774783 22.5779652502905,57.5110075378977 22.584367006355,57.4789929840942 22.6862691275745,57.3797556213022 22.7723591745184,57.390910948859 22.8511961329099,57.3784251361324 22.8697678743613,57.3844328308752 22.9189007658775,57.4218334497852 22.9485395908336,57.4058890848277 23.0078882326807,57.3669994475878 23.0110875801297,57.3549300313934 23.0247897907957,57.3541188158461 23.0327868855031,57.3438195317748 23.0358462140596,57.3372691882338 23.0484531624246))",Wilayat Bahla,ولاية بهلاء
"POLYGON ((56.001553811727 23.7843136991836,55.9583505844873 23.7867846646571,55.9556576564907 23.8254409836056,55.9191724432287 23.8209455096804,55.9145414672204 23.9153413168619,55.9017981907999 23.9516539138366,55.8697781698017 23.9256990488003,55.8508339233015 23.9551132189633,55.8206201634311 23.9551819780151,55.7954421984804 23.9616810570966,55.7810220304417 23.963387457889,55.7267899970408 24.0555296055929,55.6795353487773 24.0355849954135,55.633356567262 24.0201437480129,55.5851629548546 23.9963778022969,55.5746071827474 23.9874534331554,55.494779863629 23.9532205743413,55.4848627774221 23.9399882077393,55.498540567599 23.9237813462814,55.4996730655819 23.9076460609784,55.5123797619938 23.8948155941167,55.5245737303033 23.8772141488917,55.535175162292 23.8432848830246,55.5317855310651 23.8074073824156,55.5359026129553 23.7712348964654,55.5318400474676 23.7594902956529,55.5356219179735 23.7541190510486,55.560133672707 23.7340995631397,55.5687314577344 23.7213765933018,55.5721623127811 23.7035947689226,55.5702067175075 23.6856428589758,55.5726646075728 23.6315319101806,55.5653665548915 23.6148302189612,55.5439968711656 23.5921390142023,55.5349358637151 23.5793003920575,55.5215455712116 23.5528183397499,55.4982790791683 23.5333849299953,55.482948418695 23.5118130155712,55.4761366754871 23.4986937448198,55.4472139463608 23.4559265481205,55.4368950246114 23.4116662074322,55.4306843620394 23.3994142803459,55.4173184319815 23.3830987964139,55.531116910258 23.3356795997118,55.658966595819 23.3622815312256,55.6826707170731 23.4028437629805,55.6904625084701 23.436051834815,55.7082570786448 23.469054521229,55.7622905011625 23.4706455691061,55.8851843571015 23.5133628277196,55.975781252303 23.4981388754436,56.0109662657225 23.4792860447887,56.0334187440128 23.4988186248187,56.0534724313316 23.5338590958004,56.0325694371101 23.5530913845379,56.053603006396 23.57587050602,56.0654059990687 23.6101384860241,56.0981746644668 23.645972297091,55.9916142425238 23.7192262102091,56.001553811727 23.7843136991836))",Wilayat As Sunaynah,ولاية السنينة
"POLYGON ((56.1893392386152 24.7781721670329,56.1126963561573 24.7382043417027,56.081075900403 24.7432878292017,56.036162625135 24.8107458010023,55.9963809388683 24.8596817332573,55.9779517145884 24.8777167308196,55.9797496133316 24.8950401118457,56.0519768534689 24.87388863096,56.0418535073829 24.8887576947561,56.0407034151706 24.9089075865536,56.0633534948294 24.9478176819227,56.0415635721644 24.9468677170477,56.0458834804548 24.9681775897416,56.0300435940174 24.9733778269203,56.0066634727247 24.9945176665165,55.961023648921 25.0057278430987,55.9110902284727 24.9652994936531,55.8516160081981 24.9655265789068,55.8128681980706 24.9106974736695,55.8152486459808 24.79942305699,55.8321176110764 24.7801643045076,55.8331684634931 24.7715806819767,55.8316118417868 24.7462168319346,55.8278191451346 24.7300017139357,55.8289904574073 24.7045924820859,55.8347700230057 24.6883659862921,55.8371238996666 24.670906894145,55.7942634350144 24.6368659853362,55.8168310955927 24.6152612640302,55.7680669044049 24.5723937480196,55.7653371386759 24.5296254410144,55.7857547916398 24.4861851843026,55.8209302132916 24.4402706650151,55.827879395337 24.4099978960688,55.8346987691681 24.4100127949578,55.834424072087 24.3274339658172,55.8299604002969 24.3245630827451,55.8679265976322 24.3203618128097,55.9424360869097 24.2308079407951,55.9472184857905 24.2224983515952,55.9511854930642 24.2140720624077,55.9632886934372 24.2173807290912,55.972267213965 24.1850916300405,55.9612840580534 24.170310786512,55.975242834162 24.1461786608702,55.9956194163064 24.1254499721061,56.0149347954652 24.0898973141033,56.0132348523832 24.0877260687461,56.0178146694083 24.0674136342376,56.038114346277 24.0722049608876,56.0479139687994 24.0651352585753,56.0607040207439 24.0641682708158,56.0622363517928 24.0728920588587,56.1012159671884 24.0937699670105,56.1398343366645 24.1083155072379,56.1211765474498 24.156840154174,56.1429153523436 24.1627413515873,56.1453659820588 24.1670199635455,56.1423241792752 24.1868487347807,56.1522743185627 24.1985564538884,56.1863863386403 24.2067461890657,56.2470283805866 24.2318563247062,56.2799106579318 24.2340067593173,56.2915857356622 24.2416946448008,56.2807093972695 24.2794860850053,56.280900203305 24.3108876127464,56.3260715090555 24.3381752190403,56.342147885183 24.3758564884223,56.2807538144619 24.4242911246786,56.2242442094765 24.4278873084447,56.2188323437681 24.4872011582328,56.1969729975836 24.517662686419,56.1940279816967 24.5362507248792,56.1837813647145 24.5387829229006,56.1887000550963 24.5484193102135,56.1756850005439 24.5829685980281,56.1760236131247 24.5929498581652,56.1833670737494 24.6027228200743,56.1842378596012 24.6138157580224,56.2097985052325 24.6102247401222,56.2333464734511 24.5988863904977,56.2484956915338 24.6052082845602,56.2365390531043 24.6301300041053,56.2034970164724 24.6353560295668,56.2064895005422 24.6521272499988,56.1982916298347 24.6699479900005,56.2076150307853 24.6872456037495,56.202286165506 24.6986750552714,56.20776927219 24.7054801526812,56.2105150950118 24.7189235416316,56.2176880454103 24.7359629126459,56.2012875692826 24.749551547286,56.2017592239465 24.7601491945028,56.1902334889336 24.7699433578057,56.1893392386152 24.7781721670329))",Wilayat Mahadah,ولاية محضة
"POLYGON ((57.7183784849034 23.7693102827304,57.6670805511234 23.7759826644664,57.648074891639 23.7801014686513,57.6233041443307 23.7881205944548,57.5939428421483 23.795399748894,57.542638215424 23.8156634197434,57.5161348990359 23.8271157816073,57.5181268104177 23.812849128255,57.5386639773258 23.8030843883924,57.5257107372459 23.782162136863,57.5144974943696 23.7759008223496,57.5024876282156 23.7524071525977,57.4849876224037 23.7484042878331,57.4714990474708 23.7407654872652,57.4276118748351 23.7220477054225,57.4250709411323 23.6846540917876,57.439983535349 23.5984343054152,57.5330678986042 23.6091402681495,57.5973749106257 23.6152730935861,57.6171772165899 23.551371610473,57.6455202257619 23.5354355570249,57.6626335609093 23.609683169844,57.6901425416215 23.6508111866167,57.7015909648506 23.6936203977761,57.706691809966 23.7069414694753,57.7097746540638 23.7227570626611,57.7062917204027 23.7291241626379,57.7100203336916 23.7409557404613,57.7177334501611 23.7459156072721,57.7206573329982 23.7579930953636,57.7183784849034 23.7693102827304))",Wilayat Al Musanaah,ولاية المصنعة
"POLYGON ((57.7531923755 19.8412386672283,57.7295219109018 19.8368747901163,57.7178154461086 19.842198785119,57.7101174059157 19.8488215831795,57.6994152387587 19.8724983435129,57.6974179495321 19.8849559265303,57.6862327244957 19.9158266819629,57.6708868967224 19.9408615227175,57.6590587546202 19.94820485618,57.6307031991271 19.9518026166579,57.6090684587171 19.9585989216322,57.6029751520192 19.9795953128803,57.5958057326888 19.991450351467,57.5891253677218 19.9974140621282,57.5705401191861 19.9956608194704,57.5617988254854 20.0039396738935,57.539102582098 20.0051660987896,57.5287458907551 19.996786688145,57.5241047824191 19.9974804621947,57.4966644912685 19.9748915724979,57.4739555942643 19.9731757705178,57.4718714253564 19.9679695359023,57.4532862668901 19.964886834992,57.447617856392 19.9669095867046,57.4228216112243 19.9580174508196,57.397505336721 19.9471642867721,57.3961588160557 19.9429048861478,57.4049842306293 19.9207390298585,57.3926162757057 19.8974519376903,57.339894335995 19.8585859349464,57.3285178410388 19.7841044811833,57.3060555323464 19.7603461621647,57.2497924664554 19.5538467721999,57.1113161180224 19.3727014418215,57.0897178017582 19.3494386952711,57.0787347402994 19.3438293261446,57.0446862435819 19.335409009436,56.9864847450524 19.3185977099406,56.8635382327898 19.2792413821969,56.8031912498422 19.2567397602619,56.7494202008881 19.245426996549,56.648537834905 19.2059916058296,56.6025411008747 19.1751300734416,56.5854881638252 19.1607582717855,56.4865396656246 19.0938157204497,56.4944825157537 19.0906541909349,56.5820610094222 19.0623765655521,56.5953756307144 19.0277431016628,56.5962761385984 18.8977605347645,56.5987511151757 18.8758583969501,56.6102024668205 18.8535604132547,56.6143259136655 18.8349694649941,56.6183372888415 18.8289552317193,56.6329680366341 18.8245425769934,56.6443525575591 18.8243127110341,56.6582339708292 18.8198966243302,56.6711630370842 18.8120717143793,56.6831526076104 18.7982161021059,56.6886954373369 18.7856538729299,56.6920403287071 18.7704646208975,56.7027759237275 18.7579149129255,56.7279049354262 18.7336168010872,56.7258162668408 18.7073344536025,56.7304865372792 18.6948352731705,56.7393857038405 18.6861174159625,56.7558264453976 18.7047084062724,56.7661138703994 18.7187460906447,56.7845812395641 18.7367208887675,56.8340084111516 18.7717896874305,56.8674193489958 18.7904626456568,56.8969843058897 18.802702085464,56.9279698746064 18.8126215738773,56.9543046747487 18.8230256819021,56.9933434559928 18.8408640498685,57.0001401795441 18.8462563690659,57.0485892432088 18.8623034691224,57.0709297863688 18.8657584206747,57.107441209754 18.875737220115,57.1234972844979 18.8785346181673,57.1707370679318 18.8896430836834,57.1901636388778 18.8953970932,57.2219829609496 18.902083629673,57.2431974823268 18.9088989742341,57.286806228509 18.9191040262586,57.3134093142782 18.9234656869,57.4109655022113 18.9342507508302,57.4785795044548 18.9382606155395,57.4981200188047 18.9387130176416,57.6027190172562 18.9371250205174,57.6398356619229 18.9383292102003,57.6610438549114 18.9375036288702,57.6867872329088 18.9382799486487,57.7053085064343 18.9408391531415,57.7222531256465 18.9486419349107,57.736919800969 18.9625409530493,57.7490152223734 18.9653886345761,57.7855818134984 18.9695636931042,57.7953173882522 18.9683056786759,57.8077367463911 18.9713520005439,57.8120213593158 18.9820731853714,57.8333059864006 18.9920373592974,57.841898547943 19.0018912700048,57.8309642546434 19.0065263195175,57.821904825277 19.0165712338261,57.8150186711708 19.031238668339,57.8123761355657 19.0625549135933,57.7993673922032 19.067609158558,57.7967825121796 19.0731396453439,57.7943239063799 19.0959662047675,57.7954189290184 19.1203362347638,57.8017448960724 19.14127881149,57.8029601232576 19.1561278118313,57.792157072222 19.1697322346073,57.7765942410907 19.1675711297421,57.7624091096111 19.1830226416722,57.7535293455257 19.2086065703281,57.7510604870389 19.2243634342964,57.7441714387477 19.2321158079465,57.7407291901973 19.255173736755,57.7406546029484 19.3018645164739,57.744605509176 19.3257865971333,57.7596394162407 19.363579619718,57.7623284096419 19.3846263922064,57.7589500900606 19.409359333338,57.7532661041982 19.4281155500797,57.7484230439669 19.4326092940898,57.7475973524432 19.4450673269715,57.7404421950149 19.4495376320403,57.7317107724701 19.4664454943465,57.7263626815974 19.4691420243976,57.7197556920396 19.4942840328916,57.7017326625395 19.512284606494,57.6971189420204 19.5251626830016,57.6971086415382 19.5462383221837,57.7054414170817 19.5775027752467,57.7151738239676 19.603843957834,57.7112093705851 19.6217462083625,57.7207145068211 19.6396881642413,57.7241573952189 19.6590787567421,57.7089543676293 19.6653222797456,57.6977241939949 19.666833368531,57.6871337933922 19.6717244915377,57.6818791707675 19.6820544388132,57.677826709769 19.6993723083909,57.6769850326669 19.7119861029302,57.6839809997105 19.7381995439286,57.7014374383272 19.7629638912882,57.7371062330689 19.8006510237614,57.740524998443 19.8077843035196,57.7399304300232 19.8196236819811,57.7522910768258 19.8350865715294,57.7531923755 19.8412386672283))",Wilayat Ad Duqm,ولاية الدقم
"POLYGON ((59.0913527776265 22.7472541781927,59.0645633500111 22.7640598538002,59.047781297972 22.771610038806,59.0371374130261 22.7810804711678,59.0265462552636 22.7942166102575,59.0165985452603 22.8023435244192,58.9994445214723 22.8095603575281,58.9849324251637 22.8127526153346,58.9733634082367 22.8119424274236,58.9584895916909 22.8195846668698,58.9534225262518 22.8180530936356,58.9511835818745 22.8010939196761,58.9423418211589 22.7909121775691,58.9183450744727 22.7802124632957,58.8860903179293 22.7798809746318,58.8865129510536 22.7589204008722,58.9058120061774 22.739391154484,58.9364193046775 22.7210013925068,58.9346368834124 22.7118203971132,58.9291735128941 22.7053678973458,58.8917219938934 22.7032409712322,58.8619795249534 22.6823419822836,58.841729599172 22.6747802402113,58.8395780240146 22.6601301231717,58.8396583117527 22.6322427399342,58.8432081602316 22.6266973013434,58.8739936650135 22.599902931053,58.8847784217128 22.5860071143031,58.9009016276786 22.5580631274103,58.9025663090889 22.5469202194522,58.889617535733 22.5295289409484,58.8832565817897 22.5155068810279,58.8829370611763 22.4969844794245,58.8950488757042 22.4911516176065,58.919632659396 22.4998507053194,58.9262219812774 22.4980493133067,58.9327796940905 22.4876278075847,58.9400184361481 22.4856594436245,58.9661038543778 22.4919330389927,58.9968437811539 22.4932466999841,59.0122723234739 22.5005336368078,59.0315736550743 22.5196971210314,59.0348121129839 22.5329279527467,59.0454142858277 22.5366605509862,59.0543471702845 22.5345872373995,59.06591531823 22.5412204666424,59.084405639777 22.542568859845,59.1025486189412 22.5393845043202,59.1083267021768 22.5355751168756,59.1141053700098 22.5251219985034,59.1222644869574 22.5226186661547,59.1389875293776 22.5111830453867,59.161667340915 22.5001145713279,59.1736786927296 22.4969741318787,59.209772993222 22.4992422613091,59.2331441681103 22.5035754938877,59.2199517431622 22.5192158544764,59.2149444462081 22.5311875658368,59.2134668727311 22.5451534667415,59.2076638763575 22.5439759285805,59.1977265535305 22.5519494280398,59.1969960072709 22.5620179758383,59.2055832542139 22.5682794689524,59.205755722366 22.5869336299465,59.1930619181616 22.6045835459762,59.1799654047164 22.610423341405,59.170037231398 22.6253727384013,59.1527862499431 22.6390161007814,59.1376989123511 22.6611030236993,59.1406205141571 22.6715561222059,59.151233219355 22.6786170055577,59.1242942632743 22.7052476423795,59.1185539223589 22.7171159238787,59.1007777674698 22.7329208301466,59.0913527776265 22.7472541781927))",Wilayat Wadi Bani Khalid,ولاية وادي بني خالد
"POLYGON ((58.6499532761094 23.181007638388,58.6553744916942 23.1736400492165,58.64993211387 23.1588424558009,58.6252309641002 23.1557603258174,58.6130011825488 23.1617850176371,58.5719923704017 23.2022129480979,58.5760759733906 23.2066541371709,58.5662278435041 23.2181382244103,58.5110534888391 23.2078121959091,58.4897210743145 23.1912509287535,58.455074654626 23.2154807835916,58.4463689847575 23.2487806996584,58.4105742777666 23.2298573679404,58.4064739240594 23.223063835773,58.38338684108 23.2164818301514,58.3491418058643 23.2159816571924,58.3424045565356 23.1764488355156,58.3426395558817 23.1430943773073,58.3706095727406 23.134726495066,58.3758876507609 23.1289682572517,58.3902425127831 23.1232264317192,58.4129546179338 23.1227391722665,58.4132062422596 23.1274712554323,58.4057773447847 23.1454326342876,58.4162823274224 23.1472549325393,58.4179652119562 23.1380807717082,58.4286971866984 23.1256794074585,58.4159884598307 23.1091937338852,58.4162977432507 23.1014753389019,58.4291859175047 23.0832073518753,58.4251160816797 23.0766286251263,58.4091402519948 23.0719785082409,58.4111310665583 23.0543900266635,58.4009917258603 23.0525429579315,58.3910928129003 23.04379301979,58.3908235173287 23.035624099539,58.3781423934918 23.0278234260288,58.3760910124781 23.0143254885469,58.3846768983849 22.9998474789135,58.3760733538487 22.9847765572598,58.397511199483 22.9672641692613,58.4299074495694 22.9506889591958,58.4377564117775 22.9506586538215,58.4544506980851 22.9436877030267,58.4620456389829 22.9436562825803,58.4820313871336 22.9376049663842,58.5088615719203 22.9359161526789,58.5165129415051 22.9243125002632,58.5316457417511 22.9205885886174,58.5412728537718 22.9063005607993,58.5512153389138 22.9118234670624,58.56566065341 22.9144520434017,58.5750885516847 22.9114869127554,58.5902841619035 22.913638425248,58.5982183747665 22.9121092908446,58.6089372082733 22.9185553492451,58.6226342227425 22.9216648749318,58.6271343740227 22.9187695448594,58.6400575066581 22.9209372253533,58.6475022188731 22.9128113414371,58.6554518403269 22.9122184312225,58.6632897773327 22.9050269801826,58.6727221899272 22.9025325065768,58.6799850752812 22.9061968935971,58.6867408064557 22.9023255898273,58.6978255670053 22.9078223997699,58.709167830712 22.9062355239867,58.7233040179018 22.9085869322208,58.7377486835132 22.9152360173174,58.756265039337 22.9121244708217,58.7729697692738 22.9137472235735,58.7967811513867 22.9100819001681,58.8083995701631 22.9028250541882,58.8178715081212 22.9026763124739,58.8392093412024 22.8881876718722,58.8421195131631 22.8815302446034,58.8428701580077 22.8602890261172,58.8576323670289 22.8595890680017,58.8735971664229 22.8418764544795,58.8838302223511 22.8421868771717,58.8919602805574 22.8312000744698,58.8742916323772 22.8178049480439,58.8706335185412 22.804187398114,58.8730845940949 22.7932906772854,58.8860903179293 22.7798809746318,58.9183450744727 22.7802124632957,58.9423418211589 22.7909121775691,58.9511835818745 22.8010939196761,58.9534225262518 22.8180530936356,58.9584895916909 22.8195846668698,58.9733634082367 22.8119424274236,58.9849324251637 22.8127526153346,58.9994445214723 22.8095603575281,59.0165985452603 22.8023435244192,59.0265462552636 22.7942166102575,59.0371374130261 22.7810804711678,59.047781297972 22.771610038806,59.0645633500111 22.7640598538002,59.0913527776265 22.7472541781927,59.0899181080606 22.7528074085357,59.0909659444005 22.7752958246149,59.0874498589347 22.7852846720839,59.0749994832871 22.7962075389859,59.067280096738 22.8069276561337,59.0666613859709 22.8186085958939,59.0474775363124 22.8254050282738,59.0430700319762 22.8341503607002,59.0228794873163 22.8503455237104,59.0136686918132 22.8605868838761,59.0088044388239 22.8720485648484,58.9821420695898 22.8819715120434,58.9924621230117 22.8960851919588,58.9818551919867 22.9150894207549,58.9664441471785 22.9297611258222,58.9579629195108 22.9601451985695,58.9153821712746 22.959821037656,58.9076525564895 22.9658488218295,58.9118702581573 22.9833644344425,58.8986916559419 23.0081974511675,58.8368641958279 23.045735579718,58.8049047693354 23.0636760512512,58.7958086227328 23.1202734318818,58.7910000700562 23.125194597114,58.7919037606343 23.15277881436,58.7858179790573 23.1600310502869,58.7464969231572 23.1480524168837,58.7275880695939 23.1499790022399,58.6815602656964 23.1505744036892,58.6686140790815 23.1547878735037,58.6756257294649 23.1718062502683,58.6499532761094 23.181007638388))",Wilayat Dama Wa At Taiyin,ولاية دماء والطائيين
"POLYGON ((57.4429423167376 23.1553541340959,57.4322840535718 23.1643985881113,57.3948387209004 23.1814347312064,57.3698370217555 23.1793275261584,57.3285374807796 23.1957292645379,57.2707213717463 23.2326778043762,57.2642264609135 23.2448099945195,57.2023192742883 23.2620341670123,57.1853064160472 23.2620551664518,57.1697322393798 23.27854889679,57.1431457064386 23.2892888655115,57.1237558968639 23.2851661132575,57.0779605682882 23.2569024115974,57.0779359578782 23.2145284396679,57.0966890710622 23.2007898116578,57.1054231819287 23.1900533313597,57.115596605321 23.1883239420253,57.1201727184826 23.1774571506577,57.1332066715746 23.1714850563445,57.1385277083 23.1339107546882,57.15130461537 23.1103180353977,57.1364830571854 23.0542347628224,57.1240471750004 23.0324255196848,57.133868217636 23.0273300039486,57.1500223538638 23.0281073518141,57.1594391046784 23.0322536277856,57.1866756932885 23.0365571568731,57.2043232994765 23.0456930534614,57.2068323656364 23.0519084230132,57.2258391415713 23.0592907027261,57.227497793227 23.0793982517919,57.240914074945 23.0846407617468,57.2531973483078 23.0924724660662,57.2723047629798 23.0967141213756,57.2755310663946 23.0880526681774,57.2891911653837 23.0878774519778,57.2886851535063 23.0763366620951,57.2814620539525 23.0499244595369,57.305522226557 23.042988511844,57.3372691882338 23.0484531624246,57.3418177695608 23.0492355567763,57.3649928516505 23.0735839693801,57.3896902552256 23.0737021289662,57.4069350089254 23.0784414025226,57.4297181418011 23.1084945415168,57.4378052262602 23.1516051941218,57.4429423167376 23.1553541340959))",Wilayat Al Hamra,ولاية الحمراء
"POLYGON ((58.3760733538487 22.9847765572598,58.3846768983849 22.9998474789135,58.3760910124781 23.0143254885469,58.3781423934918 23.0278234260288,58.3908235173287 23.035624099539,58.3910928129003 23.04379301979,58.4009917258603 23.0525429579315,58.4111310665583 23.0543900266635,58.4091402519948 23.0719785082409,58.4251160816797 23.0766286251263,58.4291859175047 23.0832073518753,58.4162977432507 23.1014753389019,58.4159884598307 23.1091937338852,58.4286971866984 23.1256794074585,58.4179652119562 23.1380807717082,58.4162823274224 23.1472549325393,58.4057773447847 23.1454326342876,58.4132062422596 23.1274712554323,58.4129546179338 23.1227391722665,58.3902425127831 23.1232264317192,58.3892968043697 23.1129980902838,58.3587297362814 23.1058299505726,58.3469474898399 23.1010874746293,58.3134342280881 23.0916526960364,58.2965205679133 23.062465423235,58.2303411890025 23.0523692863411,58.2164037241019 23.052017045401,58.2071401741386 23.0452263527211,58.2012648035899 23.057314017844,58.1915319942986 23.0557095492645,58.1698539614228 23.0463262691127,58.1731934867358 23.03690684182,58.1532019979003 23.0317526076623,58.1565137868418 23.0270438975178,58.133590906604 23.0152727830984,58.1254829253822 23.0172170316306,58.0835374477787 23.0189762118738,58.050671212359 23.003650618758,58.0381539627468 22.9961158970964,58.0371092498964 22.9757761136119,58.0227409928552 22.9672022340991,58.0177028761649 22.9763317560151,58.0003491763969 22.9826034811251,57.9487417858763 22.9915292475961,57.9529666656578 22.9498597174323,57.9734289765502 22.9180215482237,57.974654914508 22.9085171004933,57.9869362174441 22.8967911833011,57.994561339742 22.8844408048127,57.9973263049985 22.8709042115709,58.011027978084 22.8638078189266,57.9948486747811 22.8428695972614,57.98876770748 22.8318062014249,57.9771333974979 22.827669082908,57.9559003499965 22.8165969614619,57.9924346854956 22.7889106780778,57.981793276584 22.7329213130798,57.9735638613173 22.7133353558484,57.9051693936022 22.6486938755621,57.90430268359 22.603321718951,57.9041180311541 22.5476842769221,57.8939798742437 22.5373745276702,57.8625786484723 22.5172629688844,57.8560468289483 22.5105368209029,57.8549500761089 22.4920868979524,57.8675006468121 22.4865379287457,57.8785060531634 22.4855646761178,57.9045408426286 22.4878387001794,57.9061786237177 22.4102653608332,57.8274075347575 22.3257127414043,57.7176454486866 22.2093141989613,57.7122144883978 22.1681812631098,57.7079918786056 22.1565414688159,57.7115601985547 22.143694602983,57.7122354734107 22.113348083222,57.6940299900165 22.1089189323367,57.6623544587289 22.0878520076207,57.6679691275807 22.0640553341978,57.7273646796641 22.0817729909505,57.7321485565712 22.0922716470253,57.7636217748654 22.0925755597166,57.7865405917639 22.0727502739145,57.8158351688434 22.0438331587693,57.8317801078301 22.0258741714211,57.8399912112635 22.00544379027,57.8618258011444 21.9581477256949,57.8823735434358 21.9079636277549,57.9197632173897 21.8589746799383,57.9437345283352 21.8285313108614,57.9670375247868 21.7724415710174,57.9675182052809 21.7373212319654,57.9392798354492 21.7240566881746,57.9439209464011 21.7003445062584,58.015357510206 21.7002713751336,58.0292212497345 21.6612086922124,58.0512449770805 21.6305955535301,58.0812254167827 21.5850850122039,58.0140813948249 21.5176959602389,58.0145450389967 21.4975344819953,58.0183138339252 21.4746774863853,58.041880705831 21.3517685337677,58.259437327468 21.4089773713887,58.2364111523592 21.4375880884629,58.2450482063561 21.453067507032,58.2656776905495 21.4550118125993,58.3574854557982 21.405577446808,58.4464065077669 21.3207835947964,58.6500242240548 21.2092389987887,58.6309980114629 21.1731215606853,58.6395427210644 21.1585215313656,58.6452329337226 21.1623014932441,58.6497504597906 21.1833056833963,58.6585153104252 21.204578716577,58.6957080005763 21.3562265299308,58.7375137006501 21.4524385866533,58.7476758227008 21.4896644423517,58.7490444530929 21.5124175651795,58.7488949047067 21.5701763461444,58.7596291065092 21.616457823968,58.7561279649038 21.6287149562157,58.7438856506011 21.6444171127965,58.7180354522144 21.668034601832,58.7088867070958 21.6858177267404,58.7049853236941 21.7126196091186,58.7095299995633 21.7425158776126,58.7163255588312 21.7600806259773,58.7280327803024 21.7990127683807,58.6914309303908 21.8401040451468,58.663448418463 21.8943650901482,58.6382493078301 21.9347779264534,58.6332896898589 21.9845666890459,58.6349931469328 22.0125510215317,58.627162210127 22.0685033509303,58.6253710632449 22.1002084916842,58.5330496789184 22.1333534559499,58.5030827707285 22.1455413559629,58.5022879082749 22.1632646297161,58.5123469298374 22.1984513556061,58.5181552632715 22.2352683770526,58.5136341545529 22.2652847912012,58.5044859247937 22.2892430839158,58.5032405217862 22.3122978730999,58.4731424346003 22.3231298443261,58.4449819339684 22.3278429074518,58.4342420881067 22.3399460162336,58.4363115682587 22.353236494051,58.4502183185346 22.3616858862897,58.4618485436933 22.3817788714014,58.5004256404748 22.4096943718055,58.5079099000624 22.4473161041588,58.4977881980113 22.4637133814487,58.4800907911352 22.4792831667778,58.4652639666239 22.5212609378503,58.4579144084094 22.5389176093836,58.4376725421565 22.5457037882681,58.4276236205336 22.5561710554946,58.4210431379664 22.5700577617672,58.3964286094309 22.5753386001599,58.3847163569436 22.5746489325737,58.3745297420688 22.5694562908617,58.3653777189842 22.5688455956304,58.358867140042 22.5729182638197,58.361431367417 22.5823089516702,58.3794078448284 22.5942165277419,58.3723627545848 22.6046876788785,58.3531837790343 22.6202565334187,58.3523298415636 22.631780837078,58.3548491910013 22.6422296463201,58.353881167675 22.6585412028102,58.3466472282369 22.675823061049,58.3463654470342 22.7011125129592,58.3514339771069 22.7101446841845,58.366084720615 22.7260919699247,58.3668716382378 22.7343655070994,58.3592720567822 22.7505622158481,58.3480450907373 22.7556691266888,58.3217517627791 22.7578500615446,58.2987238669649 22.7576032147915,58.2860712161467 22.760536735809,58.2856979410853 22.7716546049589,58.3017567588461 22.8048638031157,58.2912732238926 22.8760755458946,58.287546142367 22.8914921250943,58.293552454834 22.8913170034678,58.305720413616 22.9111118294891,58.3072899418686 22.9244089741349,58.3049550939641 22.9354491750581,58.3065854139723 22.9471703544567,58.3183499759453 22.9638798600236,58.3316191184677 22.9788873426482,58.3423127374054 22.9800687616881,58.3675501567373 22.9866421155164,58.3760733538487 22.9847765572598))",Wilayat Al Mudaybi,ولاية المضيبي
"POLYGON ((58.8510008568142 23.363473606533,58.843424876744 23.3728921273024,58.8344401879398 23.37606444084,58.8067299562262 23.3923261233206,58.7961615263127 23.4133214835574,58.784859582352 23.4234561059474,58.7780652784303 23.4644694530583,58.7797619119163 23.4740045748139,58.7762201717963 23.4847733460281,58.7628688734059 23.5017515959161,58.7616288162346 23.5122848411553,58.7199028050218 23.522132880101,58.7241680456688 23.5311680817801,58.7095662288565 23.5351438305777,58.684521695353 23.5316169847415,58.6614997679245 23.5506348580363,58.6493351304679 23.544810665642,58.6438993211718 23.5511373091729,58.6405136320433 23.5623223617888,58.6304341710067 23.5620685691155,58.6258998163293 23.5669921719722,58.6150962854277 23.569664795026,58.6064295538923 23.5812930897974,58.6017850919289 23.5945869823838,58.5989671294923 23.6167344113121,58.5919241893833 23.6180487628489,58.5850714152134 23.6251333346664,58.5711442207629 23.6227946763361,58.5778902394246 23.6133398207,58.5796017945865 23.592859512025,58.5828037693415 23.5915039547983,58.5891973948299 23.5683230908684,58.59321520152 23.5638480266928,58.5900879017391 23.5507407849228,58.592129813898 23.5416059320111,58.575522086622 23.549053599282,58.5741984274628 23.5455022213126,58.5881597371589 23.5296156981414,58.5847219754276 23.5248036403525,58.5973332833092 23.5218853266507,58.6066005917651 23.5112535927542,58.6207120472031 23.5016304521277,58.6284279137012 23.4991443029832,58.6337914657881 23.5046284533534,58.6472885230882 23.5030283020613,58.6621787776166 23.4975298828955,58.6608872950006 23.4817478351413,58.6538429551246 23.4770902163348,58.6568400938258 23.4552247486703,58.6541283952234 23.4377974934615,58.6495079369714 23.4293967135926,58.656230209715 23.4258836650048,58.6547429977717 23.4133225701908,58.6720321074424 23.4006291896654,58.6623486957117 23.38797710076,58.6655325258218 23.3793214619203,58.674774732773 23.3797713421399,58.6844763513197 23.3868050405027,58.6919014872797 23.3841083948085,58.6882046603499 23.3749218574506,58.7003403999014 23.3673541273732,58.7156719511141 23.3726704333761,58.7146580431176 23.3791607395148,58.7219419329543 23.3918132688624,58.7280476162445 23.3952766795448,58.7399596612268 23.3896158196789,58.7516019737113 23.3892826162763,58.7642001165184 23.3980603649559,58.7688223606169 23.3919467081115,58.7633051984036 23.3866293942441,58.7671407464236 23.3748831431013,58.7786089839072 23.3706851116481,58.7841861356948 23.3739175409875,58.7997365803019 23.3621403907487,58.804645081404 23.366684601093,58.8254447943019 23.3656283147251,58.8294695342696 23.3609851028518,58.8510008568142 23.363473606533))",Wilayat Muscat,ولاية مسقط
"MULTIPOLYGON (((58.6395427210644 21.1585215313656,58.6309980114629 21.1731215606853,58.6500242240548 21.2092389987887,58.4464065077669 21.3207835947964,58.3574854557982 21.405577446808,58.2656776905495 21.4550118125993,58.2450482063561 21.453067507032,58.2364111523592 21.4375880884629,58.259437327468 21.4089773713887,58.041880705831 21.3517685337677,58.070465914996 21.2024710729628,58.0387860776851 21.1401323409548,58.0140287042868 21.1143229631068,57.9910575043536 21.0496791161221,57.9946014243532 20.9407148689552,57.9851096563674 20.8977971391021,57.4665875616156 20.989135143368,57.4682687699987 20.9611358979306,57.4758836646696 20.9255703584454,57.4688672051316 20.8920358676656,57.4502551077049 20.830389544455,57.5077765667836 20.817240084704,57.5227234289762 20.8117832204638,57.5284263926757 20.7966122859438,57.5156841077731 20.772838385412,57.4328279740097 20.7752319654679,57.4108353044952 20.7287423493979,57.3658887163988 20.6974536381442,57.338163768365 20.6444713676961,57.3656944622002 20.6162720730519,57.4232271138168 20.6334595665404,57.4450548030627 20.6269101683123,57.4565040859986 20.6106439685752,57.4518225787715 20.5825132130925,57.4551874724619 20.5543612608534,57.4562756720392 20.5337922054144,57.44243704029 20.516509110218,57.4033615326527 20.5122745775466,57.4067711437722 20.4981948914322,57.3940982408966 20.4841523378482,57.3894324162231 20.4560192258095,57.3744416002119 20.4311557472657,57.3491297490045 20.4095591949979,57.3330019943814 20.3846941437157,57.3387229683337 20.3760234209214,57.3536458316756 20.3759938170831,57.3616509424294 20.3629878688884,57.3581700655025 20.3467580736534,57.348961776509 20.3348695709239,57.3718027496603 20.2882763320065,57.3889657664219 20.2698370422906,57.399231750539 20.2470820360565,57.3865456472626 20.2189660484392,57.3349347404539 20.2158246142155,57.2936258157997 20.2018261841141,57.2935710745365 20.1725990329458,57.2832083474687 20.1477186457019,57.2807517732975 20.055709923789,57.2864687898224 20.0415320276561,57.3267392886675 19.9816565419022,57.34143733598 19.9316844946072,57.3595976467853 19.9297399709134,57.3710493243599 19.9360787750025,57.3961588160557 19.9429048861478,57.397505336721 19.9471642867721,57.4228216112243 19.9580174508196,57.447617856392 19.9669095867046,57.4532862668901 19.964886834992,57.4718714253564 19.9679695359023,57.4739555942643 19.9731757705178,57.4966644912685 19.9748915724979,57.5241047824191 19.9974804621947,57.5287458907551 19.996786688145,57.539102582098 20.0051660987896,57.5617988254854 20.0039396738935,57.5705401191861 19.9956608194704,57.5891253677218 19.9974140621282,57.5958057326888 19.991450351467,57.6029751520192 19.9795953128803,57.6090684587171 19.9585989216322,57.6307031991271 19.9518026166579,57.6590587546202 19.94820485618,57.6708868967224 19.9408615227175,57.6862327244957 19.9158266819629,57.6974179495321 19.8849559265303,57.6994152387587 19.8724983435129,57.7101174059157 19.8488215831795,57.7178154461086 19.842198785119,57.7295219109018 19.8368747901163,57.7531923755 19.8412386672283,57.7676021867138 19.8716782060477,57.7710556128868 19.8842808532644,57.7687484636076 19.896783251701,57.7870021973291 19.9270721728767,57.79185968465 19.9540571889908,57.8110110410837 19.9832655226437,57.8117860291573 20.0033535127254,57.8095765278895 20.0088190984049,57.8229869053978 20.0501690155689,57.81870578641 20.0555246011287,57.8196898645665 20.0637630557897,57.832850621383 20.1039043644967,57.8315298518798 20.1143367842774,57.8344549720814 20.1249100414763,57.8193990652333 20.1382590148207,57.8145935404729 20.1695248791704,57.8241135419221 20.2010566293909,57.8466583970002 20.227122586394,57.8473612776584 20.238472543225,57.8510648877464 20.2435098187117,57.8749896613928 20.2657261853837,57.8967952174686 20.2805427231949,57.9210659159764 20.2935024518163,57.9595609521144 20.3192363525117,57.9672838939321 20.3279897457024,57.9742410343227 20.3448088121014,57.956417960596 20.3464704087582,57.9510762618448 20.350233441087,57.9428364466755 20.3668512702746,57.9438218101119 20.3860980530819,57.9485128712813 20.3969488989087,57.9571760909816 20.4079359288631,57.9761350461452 20.4224904787171,57.9937645541178 20.4318190245633,58.0277110129119 20.4450459909718,58.0479905230383 20.4495721360515,58.0550845273181 20.4577220664194,58.0621226826806 20.4584355487078,58.0672496882727 20.4691340585605,58.065715908253 20.4796704320416,58.0686479492511 20.4929155674525,58.0660718288488 20.4995082861194,58.0730069200909 20.5106038456343,58.0716750635578 20.5166774476619,58.0765780617917 20.5293742422885,58.0737195289096 20.5393620135951,58.0833404821556 20.5563803711044,58.0977859168985 20.5684887363126,58.1214285538377 20.5742279017073,58.1343673682051 20.585021432195,58.1462382211261 20.5867546601799,58.1585315729461 20.5924114659538,58.1708675004785 20.6073674314867,58.1858530348421 20.614811708599,58.2036077880961 20.6182423992486,58.2134845053654 20.6229013669763,58.2200378931507 20.620356656998,58.2287403772445 20.6048997207095,58.2578761742846 20.5953545146346,58.2736219793521 20.5807548925925,58.2806148431859 20.5785643957306,58.281667660292 20.5651970058088,58.2712316461175 20.5427533592431,58.265021733413 20.5393815122239,58.2519630807282 20.5172311096208,58.2449077107864 20.5102959216318,58.2336074752955 20.4863581752733,58.2296350516822 20.4824427339616,58.2251231383889 20.4614484681691,58.2094891378746 20.4447738432543,58.2049522402516 20.4344960784714,58.197112149064 20.4290247041441,58.2008672657854 20.4167658042952,58.1996536657333 20.4057649533119,58.2111382025998 20.3964313270264,58.224238120762 20.3948688878513,58.2728768426418 20.3747692280665,58.2823992428626 20.3684972633818,58.3018043075553 20.3758477439569,58.322576185099 20.3799377253963,58.3540916586697 20.3793323128977,58.3621209262206 20.3748203857897,58.3748559107237 20.3722563932846,58.3886312548043 20.36168109544,58.392615007414 20.3629277125146,58.4060281086597 20.3523133655039,58.4428797644952 20.3518072586773,58.4589073599579 20.3681567903253,58.4632810353568 20.3757629888963,58.474360896598 20.3828449800003,58.4755381762987 20.3912818200835,58.4831412315634 20.3930715374638,58.4917296448139 20.400347382465,58.4993519533984 20.4009708163083,58.5083266839403 20.4122489730162,58.5189084855487 20.4182142268259,58.5265187626847 20.4274818777808,58.5284952824519 20.4435379125787,58.5342857547729 20.4699919818277,58.5399914531415 20.4769855639213,58.5384098924861 20.4924427071147,58.5423094872725 20.5180005343215,58.549882240567 20.5357293038253,58.5674693796251 20.5570507152279,58.5726140565244 20.5708276332243,58.5727443639554 20.5814972872221,58.5853806749094 20.6072176506171,58.5838944515609 20.6177439435107,58.5896813687936 20.6344297060561,58.6065361984136 20.6543096464228,58.6109806924793 20.6627120882427,58.6271955348503 20.6765794622535,58.6503391356565 20.6926010395277,58.6659763317398 20.6994026613732,58.688179648076 20.713878973468,58.6984766269019 20.7286120263024,58.7126290072679 20.7426950630626,58.738375095706 20.7482290219521,58.740971136752 20.7575150693911,58.7479031540226 20.7648492715697,58.7457425224459 20.7797504075263,58.7415972087815 20.7846927699035,58.7406136076901 20.8011513447008,58.7359646785041 20.8084201288958,58.7259123806852 20.8022189855796,58.7121735019784 20.7839410028381,58.7245484885914 20.7813692258433,58.716465334108 20.7744543166719,58.7120557536146 20.7560238911687,58.7006853305689 20.7611568413215,58.6867512845523 20.7597134484256,58.6775316927059 20.7694848100023,58.6839969247462 20.7755865250894,58.6725623747306 20.7827530495816,58.6819022235166 20.7866137024328,58.6862605130953 20.7958974294828,58.6952941936269 20.8061036276537,58.6916911289159 20.8136861836936,58.7004119152288 20.8230053621103,58.7133401183873 20.8316700265423,58.7205420907845 20.8414398596778,58.7382682970212 20.8483438351332,58.7424073950408 20.855370905614,58.749640658775 20.8798919515939,58.7577431855159 20.8942293615008,58.7912631290751 20.9287180514972,58.8015451800308 20.9378584314911,58.8012955866292 20.9547615141039,58.7963849376589 20.963150830413,58.7967450851588 20.9709184766572,58.7366961758017 20.9716858835556,58.6349361204547 20.9729287941786,58.6267497461294 21.0309071231811,58.5868255477367 21.030369698721,58.6395427210644 21.1585215313656)),((58.7350003222313 20.845380929245,58.7270662589948 20.8408386397873,58.723408459802 20.8306097696775,58.7268387561825 20.8245774872807,58.7212215495759 20.8148153762556,58.7221836494102 20.8091263560361,58.7407936257224 20.8238469156026,58.7383809953219 20.8305985118622,58.739656638772 20.8450378646837,58.7350003222313 20.845380929245)),((58.1750008775651 20.5808775914434,58.163119834593 20.5813305335302,58.1637646835408 20.5722689311721,58.1702348025773 20.5660501157918,58.1759554269281 20.5698352800603,58.1750008775651 20.5808775914434)))",Wilayat Mahawt,ولاية محوت
"POLYGON ((54.6492580079343 17.2156905908809,54.6535614134464 17.2201116679904,54.6514257557516 17.2286410530679,54.6555578292206 17.2406320822791,54.6545565419886 17.2521047935051,54.6312645833698 17.2779942586386,54.6308572269503 17.3007545816364,54.6346594707051 17.3122419039691,54.6431358559315 17.3237458835882,54.6495389414065 17.3392584770749,54.655146461948 17.3399227156302,54.6595520840965 17.3514846040146,54.6529394687276 17.3591370396041,54.6442620670554 17.3553077432833,54.641589231285 17.3641216859701,54.6463263531865 17.3763301939075,54.6422515606872 17.3807635612813,54.6286940745658 17.4056757738546,54.5966548171411 17.3976313736803,54.5793335056818 17.3829066438558,54.5536707810618 17.3860486769937,54.5442848726058 17.381149654981,54.5247739590573 17.3801172376013,54.512116323299 17.3850811323603,54.4951119513884 17.370119834386,54.4741304887787 17.369855598914,54.461942388498 17.3626486907152,54.4547082668546 17.3675100181084,54.4461936134858 17.3667716361368,54.4384980886349 17.3542889647882,54.4291013225838 17.3541683256386,54.4179288791555 17.3403809539426,54.41683514964 17.3248343696144,54.4121165409057 17.3184764925348,54.3932619605621 17.3228496310698,54.3841703201751 17.3321762578768,54.3710128745194 17.335362096216,54.3538137863553 17.3460495929237,54.3547346923736 17.3580254547748,54.3498397339335 17.3640473673101,54.328029899255 17.3608184555843,54.3306068324161 17.348889417749,54.3208991169093 17.3401543011274,54.3101471152306 17.3431582368418,54.3049921496272 17.3370022500973,54.3049482995579 17.3250383638969,54.2849693200102 17.3165830499782,54.2897385130626 17.3042646999342,54.2854421061579 17.2952907445055,54.2891411883231 17.2894447492353,54.2904173529812 17.2770173923312,54.2853202980322 17.2683059316176,54.2890175489326 17.2616256020981,54.2989925146391 17.2604674106444,54.3149205979886 17.2657249271423,54.3228112012221 17.2487549340234,54.3209066202708 17.2327582820497,54.3161534078258 17.2319024834728,54.3075570833379 17.246014250337,54.2962410048205 17.2490115069487,54.2941323834261 17.2249116276991,54.2796950193499 17.2126769404264,54.281410374647 17.2045554003689,54.2956604217455 17.2020846990975,54.3051923093605 17.1816712793552,54.2754722424394 17.1397571703852,54.2678642142944 17.1311820699552,54.269797372398 17.1223002168863,54.2651791601233 17.1115737047415,54.2573261263924 17.1075889511152,54.2544756250448 17.1009867482311,54.2432687084464 17.098111528152,54.2335184422624 17.090759979966,54.2387275312855 17.0717610220964,54.2491898469013 17.0532716302036,54.2681718308247 17.0506532870678,54.2749356449547 17.0543152171232,54.2986087029291 17.0531505822188,54.3205983168218 17.0620596955423,54.3316265609454 17.0642248219803,54.3420296783292 17.0611297539931,54.3394810429385 17.0532865288308,54.341918296573 17.0316897681505,54.4087079482171 17.0335071325859,54.4368306782718 17.0306943360123,54.4305192393024 17.0380261217018,54.4260397039182 17.0489804314376,54.4240594077781 17.067380196003,54.4278031890652 17.0770172446557,54.4385613030032 17.0761053530663,54.4400437852001 17.0857871846345,54.4476674413374 17.0871074070476,54.4532094511681 17.0939769787428,54.4587811007486 17.113114536144,54.4718020132633 17.1372756131967,54.4732587900349 17.1461746557213,54.4718253515884 17.1625849009286,54.4897827262511 17.1618252247125,54.4974933923401 17.1644889165798,54.5029783021952 17.1718628080508,54.5134483907022 17.1726661391802,54.5366134979891 17.1832032873037,54.5430090614854 17.1819591914119,54.5516870325872 17.1876667960139,54.5604463440145 17.177450088391,54.568203943219 17.1929357136393,54.5800318932545 17.1976529908274,54.5845908524128 17.2082849539881,54.5922609891093 17.1991662781376,54.6044756221806 17.1995661880842,54.60655628544 17.2123893043833,54.6139702461963 17.2077804326205,54.6329423612385 17.2072785895411,54.6384666407179 17.2177970511788,54.6492580079343 17.2156905908809))",Wilayat Taqah,ولاية طاقة
"POLYGON ((55.2576537967518 17.5856522039584,55.2418539779035 17.5848660907932,55.2187004461355 17.589924193437,55.2132518976959 17.5775529702305,55.1821072379549 17.5616154557882,55.1719596732682 17.5499794315076,55.16219229904 17.5514351687196,55.1426497320786 17.5480351644398,55.1263580088269 17.5391289541604,55.1079086198521 17.5410135888607,55.0894498591354 17.5331815747766,55.0847404972227 17.5261250230731,55.0615707899427 17.5044342055981,55.0499928227394 17.5001421873469,55.0405836449177 17.492827376509,55.0282854267199 17.4914972445805,55.0167092383805 17.4872034388091,55.0083867803474 17.4793549117274,54.9935570746075 17.4742525182301,54.9758312914071 17.4590857061596,54.9494360474582 17.4662088113574,54.9443748511466 17.4752032941355,54.9378658453956 17.4769788537789,54.9309941352328 17.4700255733846,54.9234010088732 17.481567793684,54.9139983254251 17.4815359122032,54.9082121119103 17.4881388811761,54.8912135954757 17.4972212771719,54.8760228906223 17.5018541033096,54.8774649277586 17.5231592249447,54.8742084979148 17.5272009023758,54.8608248443965 17.5273708362937,54.8539458966492 17.5451947757681,54.8430943917676 17.5432825435078,54.8289854636611 17.5449418994004,54.828259917625 17.549350298537,54.8137890337966 17.5505257546532,54.7895577567849 17.5424551125644,54.7302275143275 17.5496666469323,54.713948251636 17.5509325389987,54.6893776516345 17.5297494037554,54.6756211172857 17.5391476333843,54.6705630002873 17.5350143676777,54.6636993198256 17.5290203946992,54.6470575913315 17.532244669684,54.6427009136416 17.5431315607886,54.6358229520044 17.5468602465519,54.6275164172852 17.5389972989193,54.6271740840006 17.5268656902998,54.6152720109076 17.5070237924173,54.6178304595637 17.4903825002186,54.6127862565292 17.4794511307398,54.6193088951347 17.4703984901142,54.6193204068271 17.4631115048723,54.6258353976599 17.4584314192187,54.6254933861438 17.4458210235288,54.6305834086636 17.4266339827413,54.639292977886 17.4029031289065,54.6286940745658 17.4056757738546,54.6422515606872 17.3807635612813,54.6463263531865 17.3763301939075,54.641589231285 17.3641216859701,54.6442620670554 17.3553077432833,54.6529394687276 17.3591370396041,54.6595520840965 17.3514846040146,54.655146461948 17.3399227156302,54.6495389414065 17.3392584770749,54.6431358559315 17.3237458835882,54.6346594707051 17.3122419039691,54.6308572269503 17.3007545816364,54.6312645833698 17.2779942586386,54.6545565419886 17.2521047935051,54.6555578292206 17.2406320822791,54.6514257557516 17.2286410530679,54.6535614134464 17.2201116679904,54.6492580079343 17.2156905908809,54.6639259200827 17.2139542170614,54.6683338186417 17.2075037068209,54.6920657187022 17.2039345318292,54.7209930075119 17.1877993205202,54.7324913959998 17.1840953808622,54.7489952200119 17.1746933925409,54.7599050168269 17.1656761545955,54.7956538492785 17.1544725507919,54.8034141993748 17.1532087978056,54.8110913501748 17.1569057177508,54.8222409103796 17.1566886240163,54.8243435040524 17.1451692292661,54.8202302286665 17.1323545908742,54.8396917895009 17.1226969741735,54.8422950951509 17.1108646351996,54.8422482581324 17.0792370857004,54.8539180756724 17.0670929955623,54.8590329679966 17.057722514217,54.8604608292539 17.0470564242474,54.8684805600494 17.0310142313611,54.871454819671 17.0182698075338,54.8683463626252 17.0044144825633,54.8627470199481 16.999119875721,54.8494664825895 16.9993988875312,54.842870194602 16.9953156997091,54.8484722407514 16.9815723843413,54.8583032294457 16.9641125038756,54.8705216875916 16.9605536036772,54.8780607688676 16.9685542085286,54.8872935828739 16.965070181751,54.9046173653128 16.9677367927541,54.9115327114852 16.978634523788,54.9132559182874 16.9915128678956,54.9245681052414 16.9829970172139,54.9270606765633 16.9771058392986,54.9374800819845 16.9781522795792,54.9431348761608 16.989404550703,54.9566041299611 16.9871063792394,54.9687071347481 16.9905488450478,54.9838246858194 17.0018650338939,54.9912952483953 17.0217321038115,55.0091066419186 17.0207245463242,55.0210778771206 17.0140015978391,55.0258317822179 17.0064903542754,55.0340448883712 17.0165752372927,55.040202645379 17.0190225026572,55.0578652561881 17.0336517644544,55.0733434422461 17.0397311026512,55.0761787248189 17.0460323840453,55.0841641438199 17.0475726910844,55.0856492191474 17.057464500066,55.1003142276493 17.0671469402822,55.1204855951253 17.0892483440262,55.1263420089638 17.1039203386114,55.1354765350789 17.1111656494816,55.1420197546576 17.1263300460855,55.1609123178852 17.13670360446,55.1869938379202 17.141628253755,55.1928026276863 17.1484559044349,55.1930386995703 17.1625412417494,55.2050559426655 17.1776127245099,55.2052428771187 17.1825845666504,55.2142529969343 17.1938122839871,55.229085100833 17.199963854086,55.237265486323 17.2111683276418,55.246481766072 17.2169442503283,55.2531960394448 17.2310193028268,55.2628219930137 17.2442182337926,55.2566031392971 17.2471293007642,55.2419560305073 17.2673232427739,55.2424861695284 17.279661721161,55.2493734051413 17.2934280827399,55.2620201812738 17.2982118548116,55.2672489083493 17.3196280149464,55.2782207983127 17.330277661997,55.2800744361808 17.3485460603386,55.2941683070842 17.3590546710897,55.2921152927645 17.3681001516131,55.2988586354937 17.3787940794055,55.2968794723534 17.3902415130038,55.3013636115211 17.3951026422321,55.2956846618086 17.4080997782735,55.2847604964888 17.4247254751284,55.2818704018572 17.4367460270908,55.2714467794306 17.4493972281691,55.2608168811478 17.4473889528073,55.2428342315512 17.4530325110386,55.2308782488815 17.4722591765228,55.2302633484519 17.4976994102624,55.225544475829 17.5024472463421,55.2236623447375 17.5180641004792,55.2274294746286 17.5374281503705,55.2388394119865 17.5634031599361,55.2576537967518 17.5856522039584))",Wilayat Sadah,ولاية سدح
"POLYGON ((54.7725551691783 18.4590161358455,54.0462645146381 19.2764483805776,53.7610341920431 19.5941902700002,53.6289915058907 19.5503381151519,52.6178205315456 19.2107400398903,53.0059225643277 18.4250246465511,53.1786469516003 18.158622745698,53.1716091983395 18.1554783499491,53.1485757690599 18.1231586341157,53.1352993254534 18.1128974098772,53.1061469315797 18.1116850638238,53.0888721914108 18.0757293811523,53.0815653478731 18.0518442107512,53.0816047759337 18.0206123531318,53.0804220551131 17.9953940255254,53.0608885107734 17.983337389818,53.056238075992 17.9674185133832,53.0586941083733 17.9449813861158,53.035491824974 17.903043171822,53.0373745787168 17.8380991038042,53.0601359284356 17.8179966629723,53.0586426459524 17.7726459486622,53.0495145332738 17.7422752050237,53.0351258915459 17.7418967033466,53.0131563609995 17.7322392695085,53.0200898319925 17.7196256607608,53.0419947628093 17.7147352383439,53.043965042266 17.6978987426785,53.0728240445654 17.6895849028656,53.0832410540031 17.6882894267513,53.0934330603625 17.6661588143249,53.0989887983042 17.6347072840721,53.0918866602642 17.6172407249011,53.0921941195988 17.5960836239516,53.0877830999771 17.5920796728692,53.1052157204988 17.549854873121,53.13873965963 17.510436914113,53.1866057968622 17.468078433119,53.187019694369 17.4482122210308,53.1587031772243 17.4374010060192,53.1438801057085 17.4219681978746,53.1359852959352 17.4072750634862,53.1362528475868 17.3945577211089,53.1409096324381 17.3831370235225,53.1493623994071 17.3711835447282,53.1570063390376 17.3676958217968,53.1708558277822 17.3691737253947,53.1757628030639 17.3759322643165,53.1883792625443 17.3827702062217,53.2273317908702 17.4086275548016,53.2342443948302 17.4164277223108,53.2429900362876 17.420834214738,53.2574763253113 17.4223188986933,53.2838528144845 17.4288722751175,53.306726428933 17.4214210060459,53.3196250222885 17.4077232793871,53.323321433409 17.3934881805661,53.3155784609245 17.3829575262929,53.3147141446429 17.3682020232057,53.3110833691642 17.3647799505993,53.2938060606769 17.3626262675592,53.2815193150336 17.3529607395593,53.2394022643881 17.3287895552054,53.2193630663332 17.3113276673099,53.2059146222433 17.2904733095492,53.2063649533133 17.2778942718223,53.2184375366874 17.2640510229503,53.2292522489713 17.2594074161648,53.2405985698011 17.2596202845928,53.2675822623849 17.2661831105396,53.2819112423453 17.274932108825,53.2984191223436 17.2994913896907,53.3127394005391 17.313786146466,53.3408457299294 17.3244926117212,53.3624074228069 17.3188261770836,53.3708914925266 17.3044368875603,53.3680954988911 17.2862070609766,53.3464939694612 17.2688042007644,53.3414617118442 17.2614843988831,53.337335979827 17.2468662055182,53.3407627049203 17.2329916318333,53.3555221635339 17.2199285567752,53.3745260445819 17.2154242283351,53.4133356390444 17.2191757117935,53.4899248996613 17.2140640098801,53.5447132433727 17.2190256413875,53.557344373748 17.2180300745752,53.5987859585823 17.221570996105,53.6424681290096 17.2188627725109,53.6613940146887 17.2185716417436,53.6673934811591 17.2316886011198,53.6615280342989 17.2563388438214,53.6601148113017 17.2778076253579,53.6665573915732 17.3070222488302,53.67567233767 17.3129293909364,53.677365214105 17.3215215551348,53.6865978021781 17.3266935017429,53.6883963420857 17.3403164421637,53.6977275412071 17.3526039512653,53.7025186175328 17.354576456834,53.7185054882494 17.3492068436696,53.7267176694247 17.349467896199,53.7396339737321 17.338079169475,53.7457914677733 17.3396836250074,53.7527392339117 17.3482844323302,53.7609621740432 17.3444943797938,53.7592646654137 17.336270099235,53.7637234827456 17.3303876607074,53.7737665960961 17.3295444578193,53.77947815147 17.3215772408585,53.7733313491702 17.3129789409858,53.7712907404443 17.3029132324317,53.7820264258755 17.2969168296695,53.7944554346466 17.3000026038715,53.8114642170068 17.2942581841208,53.8278920744539 17.2958741705483,53.8313208638521 17.2891293263611,53.8455789845279 17.2897593144402,53.8623421859599 17.2975089057648,53.8705377684425 17.2942296291276,53.8744135739319 17.2727360713367,53.8803758162338 17.2536350872251,53.8931164257033 17.2489713631281,53.9106632832009 17.2516800730667,53.9304797601486 17.2657838110179,53.9345902430802 17.26014169033,53.9475952578047 17.2576944208784,53.9615151154785 17.2591752035256,53.9675599893085 17.2562329027845,53.9862695321431 17.2585731475514,54.0006415945691 17.264223822301,54.0207219691201 17.2676661232327,54.0313343444464 17.2654599613999,54.0432006018716 17.2668111685027,54.0489037260466 17.2733172360524,54.0580324258778 17.277122874612,54.0640824092207 17.2902556859941,54.0732120963866 17.293201865658,54.0824586922949 17.3037567839174,54.0902192418542 17.3033888145211,54.0931781092977 17.3104768093685,54.1030021857853 17.3058416351551,54.1071124841193 17.311119086235,54.1646061086162 17.3120158811322,54.1773640470004 17.3190185200815,54.1937907210464 17.3316071753453,54.2034319109691 17.3314127519617,54.2094739785077 17.3385032888999,54.227206944813 17.3524606353065,54.2426953111585 17.3692297386697,54.2684013412137 17.4048525518844,54.2806217314327 17.4402893815305,54.2915698093844 17.4605929446169,54.2973239322992 17.4772265719369,54.2935888165975 17.526841438044,54.2868143911518 17.548473099296,54.3514599310961 17.5307456863914,54.4228278168332 17.5355249610325,54.5048805631248 17.5535734989527,54.5661347306943 17.5894300857515,54.616812259086 17.6380342415251,54.5406116650914 17.6977655254461,54.5136290703897 17.7114747897224,54.4927119860155 17.7323475810809,54.4665227647879 17.7452061304034,54.4527968266192 17.7420960712777,54.3771468595672 17.6839234991748,54.3575687619713 17.6631371277314,54.3348082841046 17.6511022765099,54.3105659823764 17.6361129677918,54.2816107799332 17.6298519302902,54.2540978128588 17.6294706372033,54.218920878316 17.6304434171166,54.182170544389 17.6343190708565,54.1590375324419 17.6471793673281,54.1404409407861 17.6630340507496,54.1463009726096 17.6792429638513,54.1613813982375 17.6926535952775,54.1978251162553 17.7093010271851,54.2268329707826 17.712644595219,54.2587003695491 17.7292171836693,54.2832111020304 17.7467608756346,54.2856922895049 17.7612170503241,54.3004883205712 17.798696338944,54.3245963666066 17.8239491879316,54.4425749843145 17.9222907886722,54.5242820891021 17.989734493238,54.5538176644689 17.9890229688734,54.5802941117621 17.9805266607265,54.6017358753032 17.9543064583193,54.6139155066845 17.9304922156928,54.635496252286 17.8929169780122,54.6552537792696 17.8931559631988,54.6721303133851 17.9122784555583,54.6994459430645 18.0412603029575,54.7001403539192 18.0891991888459,54.6586754414776 18.1328456198315,54.6389419024359 18.1288206782273,54.585230697132 18.1016682316831,54.5453086786816 18.0915861209749,54.5472283165309 18.1069087014806,54.5465277832101 18.1507048736303,54.5563120785597 18.1594266510923,54.5536135974793 18.196153982824,54.5677151275365 18.2281005346707,54.624220367658 18.2950962935969,54.643518501198 18.3220537015553,54.6595662044005 18.3411117448775,54.7225730898391 18.4003292053433,54.7557209310514 18.4350149264513,54.7633703001456 18.4553294145187,54.7725551691783 18.4590161358455))",Wilayat Thumrayt,ولاية ثمريت
"MULTIPOLYGON (((56.3536691272746 17.9210449091626,56.3450819376393 17.9329781413001,56.0237167595048 18.4326668676184,56.0149679382374 18.4462205857403,55.9670214285953 18.4419598478503,55.951247638415 18.4446293580058,55.946630604823 18.4528472131174,55.9445406989223 18.4698909425214,55.958120296298 18.4738509281263,55.9694533515313 18.4725950319863,55.9946283204056 18.4777204910562,56.0003783363524 18.4841592644063,55.9979481760327 18.5073924624753,55.9858954350691 18.5152453306629,55.9684209435662 18.5182865053955,55.9270805938945 18.5090223145744,55.8828463880479 18.4969635441073,55.868387156205 18.4903662564688,55.8515155336813 18.4920628717873,55.8413951844763 18.4897889958427,55.7663842739647 18.5989966326859,55.8565817421901 18.6911301010414,55.8402280132996 18.7163673047502,55.6891378079147 18.9490818683714,55.3579352899718 18.9313324723516,55.2287822075882 18.9256701840039,55.1166023246808 18.9219061973567,55.0781669397002 18.8987065213805,55.0661983983014 18.8784710557405,55.0277972884834 18.8563973757166,55.0001456251945 18.8443599826372,54.9975942516966 18.8160217276074,54.9921031628097 18.8002185110969,54.9759114607706 18.7766414513007,54.9518388834975 18.7214068071312,54.9546843242214 18.6997928398827,54.9086953521663 18.6596602408353,54.8784559444168 18.6124631062867,54.8560576436228 18.5969198042189,54.81118371301 18.5567518641076,54.808825292255 18.5374924935908,54.7853783843904 18.5219604618106,54.7872110223373 18.5003677105381,54.7824422325126 18.4629840636509,54.7725551691783 18.4590161358455,54.7633703001456 18.4553294145187,54.7557209310514 18.4350149264513,54.7225730898391 18.4003292053433,54.6595662044005 18.3411117448775,54.643518501198 18.3220537015553,54.624220367658 18.2950962935969,54.5677151275365 18.2281005346707,54.5536135974793 18.196153982824,54.5563120785597 18.1594266510923,54.5465277832101 18.1507048736303,54.5472283165309 18.1069087014806,54.5453086786816 18.0915861209749,54.585230697132 18.1016682316831,54.6389419024359 18.1288206782273,54.6586754414776 18.1328456198315,54.7001403539192 18.0891991888459,54.6994459430645 18.0412603029575,54.6721303133851 17.9122784555583,54.6552537792696 17.8931559631988,54.635496252286 17.8929169780122,54.6139155066845 17.9304922156928,54.6017358753032 17.9543064583193,54.5802941117621 17.9805266607265,54.5538176644689 17.9890229688734,54.5242820891021 17.989734493238,54.4425749843145 17.9222907886722,54.3245963666066 17.8239491879316,54.3004883205712 17.798696338944,54.2856922895049 17.7612170503241,54.2832111020304 17.7467608756346,54.2587003695491 17.7292171836693,54.2268329707826 17.712644595219,54.1978251162553 17.7093010271851,54.1613813982375 17.6926535952775,54.1463009726096 17.6792429638513,54.1404409407861 17.6630340507496,54.1590375324419 17.6471793673281,54.182170544389 17.6343190708565,54.218920878316 17.6304434171166,54.2540978128588 17.6294706372033,54.2816107799332 17.6298519302902,54.3105659823764 17.6361129677918,54.3348082841046 17.6511022765099,54.3575687619713 17.6631371277314,54.3771468595672 17.6839234991748,54.4527968266192 17.7420960712777,54.4665227647879 17.7452061304034,54.4927119860155 17.7323475810809,54.5136290703897 17.7114747897224,54.5406116650914 17.6977655254461,54.616812259086 17.6380342415251,54.6520646719631 17.596488477638,54.6645766868259 17.5746421919644,54.6705630002873 17.5350143676777,54.6756211172857 17.5391476333843,54.6893776516345 17.5297494037554,54.713948251636 17.5509325389987,54.7302275143275 17.5496666469323,54.7895577567849 17.5424551125644,54.8137890337966 17.5505257546532,54.828259917625 17.549350298537,54.8289854636611 17.5449418994004,54.8430943917676 17.5432825435078,54.8539458966492 17.5451947757681,54.8608248443965 17.5273708362937,54.8742084979148 17.5272009023758,54.8774649277586 17.5231592249447,54.8760228906223 17.5018541033096,54.8912135954757 17.4972212771719,54.9082121119103 17.4881388811761,54.9139983254251 17.4815359122032,54.9234010088732 17.481567793684,54.9309941352328 17.4700255733846,54.9378658453956 17.4769788537789,54.9443748511466 17.4752032941355,54.9494360474582 17.4662088113574,54.9758312914071 17.4590857061596,54.9935570746075 17.4742525182301,55.0083867803474 17.4793549117274,55.0167092383805 17.4872034388091,55.0282854267199 17.4914972445805,55.0405836449177 17.492827376509,55.0499928227394 17.5001421873469,55.0615707899427 17.5044342055981,55.0847404972227 17.5261250230731,55.0894498591354 17.5331815747766,55.1079086198521 17.5410135888607,55.1263580088269 17.5391289541604,55.1426497320786 17.5480351644398,55.16219229904 17.5514351687196,55.1719596732682 17.5499794315076,55.1821072379549 17.5616154557882,55.2132518976959 17.5775529702305,55.2187004461355 17.589924193437,55.2418539779035 17.5848660907932,55.2576537967518 17.5856522039584,55.2582231837607 17.5971713095387,55.2634651579642 17.6039670454203,55.2904270144251 17.6221991206133,55.3020876885809 17.6285412344622,55.3027596139775 17.6351555172803,55.3146810454494 17.6443771089521,55.3191930442878 17.6512444216225,55.3423949796589 17.6607513009262,55.3547670316916 17.668418085302,55.3557886854286 17.6723865989445,55.3767550394176 17.6806410353692,55.376280027167 17.688168581183,55.3846296027763 17.7033003035878,55.3796501399401 17.7107489813762,55.3805985234327 17.7291584884501,55.3927459906174 17.7487590785912,55.4014456484979 17.7516494196993,55.4145700556779 17.7614776235545,55.4172031236078 17.7722777626167,55.4132268587783 17.7816735344084,55.4207378531702 17.7990924659182,55.418985914705 17.8065680338759,55.4265802769938 17.8181423136188,55.4436018622409 17.8247699042857,55.4868003159522 17.8466832245862,55.5261692040616 17.8608213780563,55.5511769580163 17.868678400489,55.5879780614381 17.8781904656279,55.6295007451505 17.8866682270295,55.6656817306332 17.8915205137136,55.7188752824626 17.896217807619,55.7295864987741 17.8997365597402,55.7497636712989 17.9020812429932,55.7853138445796 17.9026892722684,55.8299504528105 17.900411949937,55.8402203871937 17.898922390243,55.8526282185938 17.9011399966183,55.8670810790575 17.896460861368,55.8912364262054 17.8938886996427,55.9109188573212 17.896689524486,55.9302763210363 17.9039228584751,55.9445059827892 17.9166699441595,55.9737148308823 17.9261631328828,55.9781726244917 17.9302535008102,56.0125967943015 17.9285583490238,56.0191185160518 17.930672274541,56.0631572060456 17.9275929819009,56.0997101715962 17.921134374488,56.1091921772538 17.9216343540665,56.1143336774073 17.9269609624929,56.1459092333772 17.9276717015779,56.1555181886774 17.9312881646632,56.1647497710059 17.939716950631,56.2301631475635 17.9382422236457,56.2780641844755 17.9326467409871,56.2798677097877 17.9282307157927,56.2918253166988 17.926817506486,56.3052654734783 17.9212639533638,56.322386782683 17.9179469614025,56.3441213893985 17.9172595697635,56.3536691272746 17.9210449091626)),((56.0506814740479 17.5539438481717,56.0331000075304 17.5383936362707,56.0137136380429 17.5295157725642,55.9930561890261 17.5280320191962,55.9767688073508 17.5187671290051,55.9637861572693 17.5146673088901,55.9638474412064 17.495369231756,55.9819867905818 17.4903573393557,55.9905756714366 17.4847493762552,56.0090824992824 17.4840201655851,56.0122880455036 17.4798798163447,56.0330277784928 17.479844923469,56.0569224962928 17.4883459742374,56.0707550195433 17.4959026335821,56.0883825388335 17.5009327258798,56.0936062957812 17.5128034127384,56.0825066514978 17.51087133778,56.0625039311923 17.5154019600092,56.0557286868234 17.5344819482888,56.0560179199584 17.5458882192447,56.0506814740479 17.5539438481717)),((55.8488926989085 17.5086629809965,55.8254012920493 17.4933004785647,55.8267881093837 17.4858651262667,55.8438843987827 17.4834958224069,55.8508204507959 17.4881350729806,55.8606312353626 17.476691184247,55.8738270379555 17.4769121180261,55.882030017335 17.485601852728,55.8798482788675 17.4953660782961,55.8700214221094 17.4951375615072,55.8617102543043 17.5026319983377,55.8488926989085 17.5086629809965)),((56.3402943274425 17.507980934328,56.3329637704546 17.5081711001091,56.3237214955574 17.4985114783848,56.3381892543835 17.4957085450355,56.3434944674518 17.4911706901852,56.3527366101663 17.4966637408486,56.3477347133921 17.5061322731032,56.3402943274425 17.507980934328)),((55.6037409091094 17.4848814459779,55.5946890776887 17.4810266572109,55.5962028704063 17.4698519546974,55.6051908435539 17.4720580895882,55.6096876560508 17.479155334557,55.6037409091094 17.4848814459779)))",Wilayat Shalim Wa Juzor Al Hallaniyat,ولاية شليم وجزر الحلانيات
"POLYGON ((54.6492580079343 17.2156905908809,54.6384666407179 17.2177970511788,54.6329423612385 17.2072785895411,54.6139702461963 17.2077804326205,54.60655628544 17.2123893043833,54.6044756221806 17.1995661880842,54.5922609891093 17.1991662781376,54.5845908524128 17.2082849539881,54.5800318932545 17.1976529908274,54.568203943219 17.1929357136393,54.5604463440145 17.177450088391,54.5516870325872 17.1876667960139,54.5430090614854 17.1819591914119,54.5366134979891 17.1832032873037,54.5134483907022 17.1726661391802,54.5029783021952 17.1718628080508,54.4974933923401 17.1644889165798,54.4897827262511 17.1618252247125,54.4718253515884 17.1625849009286,54.4732587900349 17.1461746557213,54.4718020132633 17.1372756131967,54.4587811007486 17.113114536144,54.4532094511681 17.0939769787428,54.4476674413374 17.0871074070476,54.4400437852001 17.0857871846345,54.4385613030032 17.0761053530663,54.4278031890652 17.0770172446557,54.4240594077781 17.067380196003,54.4260397039182 17.0489804314376,54.4305192393024 17.0380261217018,54.4368306782718 17.0306943360123,54.4878389942082 17.0341027047856,54.5011927559823 17.0328856821128,54.5263443840114 17.0335809189907,54.5440567048216 17.0306564385001,54.558882503686 17.0316617496197,54.5682152370345 17.0290098117324,54.5818764805116 17.0298329294059,54.6379005337221 17.0252018663163,54.6589451517591 17.0209857552779,54.6750208705317 17.0159133222281,54.6843353494248 17.0092798610889,54.6910379012648 16.9915784661842,54.6838112393872 16.9821116837798,54.6846764393607 16.9770679326182,54.6963204824726 16.9741824898035,54.6967842902666 16.9670062901429,54.7111712340659 16.9687184883702,54.7317532417435 16.9592826632907,54.7400193016639 16.9522434425848,54.7562309844713 16.9608369317557,54.765669302256 16.9521782374266,54.7773543524283 16.9554266501039,54.7838582084266 16.9537277456777,54.7993394578199 16.9414567781079,54.8173413144276 16.9499410660472,54.8151224598886 16.9559408103261,54.828916463354 16.9628783608085,54.8583032294457 16.9641125038756,54.8484722407514 16.9815723843413,54.842870194602 16.9953156997091,54.8494664825895 16.9993988875312,54.8627470199481 16.999119875721,54.8683463626252 17.0044144825633,54.871454819671 17.0182698075338,54.8684805600494 17.0310142313611,54.8604608292539 17.0470564242474,54.8590329679966 17.057722514217,54.8539180756724 17.0670929955623,54.8422482581324 17.0792370857004,54.8422950951509 17.1108646351996,54.8396917895009 17.1226969741735,54.8202302286665 17.1323545908742,54.8243435040524 17.1451692292661,54.8222409103796 17.1566886240163,54.8110913501748 17.1569057177508,54.8034141993748 17.1532087978056,54.7956538492785 17.1544725507919,54.7599050168269 17.1656761545955,54.7489952200119 17.1746933925409,54.7324913959998 17.1840953808622,54.7209930075119 17.1877993205202,54.6920657187022 17.2039345318292,54.6683338186417 17.2075037068209,54.6639259200827 17.2139542170614,54.6492580079343 17.2156905908809))",Wilayat Mirbat,ولاية مرباط
"POLYGON ((54.6705630002873 17.5350143676777,54.6645766868259 17.5746421919644,54.6520646719631 17.596488477638,54.616812259086 17.6380342415251,54.5661347306943 17.5894300857515,54.5048805631248 17.5535734989527,54.4228278168332 17.5355249610325,54.3514599310961 17.5307456863914,54.2868143911518 17.548473099296,54.2935888165975 17.526841438044,54.2973239322992 17.4772265719369,54.2915698093844 17.4605929446169,54.2806217314327 17.4402893815305,54.2684013412137 17.4048525518844,54.2426953111585 17.3692297386697,54.227206944813 17.3524606353065,54.2094739785077 17.3385032888999,54.2034319109691 17.3314127519617,54.1937907210464 17.3316071753453,54.1773640470004 17.3190185200815,54.1646061086162 17.3120158811322,54.1071124841193 17.311119086235,54.1030021857853 17.3058416351551,54.0931781092977 17.3104768093685,54.0902192418542 17.3033888145211,54.0824586922949 17.3037567839174,54.0732120963866 17.293201865658,54.0640824092207 17.2902556859941,54.0580324258778 17.277122874612,54.0489037260466 17.2733172360524,54.0432006018716 17.2668111685027,54.0313343444464 17.2654599613999,54.0207219691201 17.2676661232327,54.0006415945691 17.264223822301,53.9862695321431 17.2585731475514,53.9675599893085 17.2562329027845,53.9615151154785 17.2591752035256,53.9475952578047 17.2576944208784,53.9345902430802 17.26014169033,53.9304797601486 17.2657838110179,53.9106632832009 17.2516800730667,53.8931164257033 17.2489713631281,53.8803758162338 17.2536350872251,53.8744135739319 17.2727360713367,53.8705377684425 17.2942296291276,53.8623421859599 17.2975089057648,53.8455789845279 17.2897593144402,53.8313208638521 17.2891293263611,53.8278920744539 17.2958741705483,53.8114642170068 17.2942581841208,53.7944554346466 17.3000026038715,53.7820264258755 17.2969168296695,53.7712907404443 17.3029132324317,53.7733313491702 17.3129789409858,53.77947815147 17.3215772408585,53.7737665960961 17.3295444578193,53.7637234827456 17.3303876607074,53.7592646654137 17.336270099235,53.7609621740432 17.3444943797938,53.7527392339117 17.3482844323302,53.7457914677733 17.3396836250074,53.7396339737321 17.338079169475,53.7267176694247 17.349467896199,53.7185054882494 17.3492068436696,53.7025186175328 17.354576456834,53.6977275412071 17.3526039512653,53.6883963420857 17.3403164421637,53.6865978021781 17.3266935017429,53.677365214105 17.3215215551348,53.67567233767 17.3129293909364,53.6665573915732 17.3070222488302,53.6601148113017 17.2778076253579,53.6615280342989 17.2563388438214,53.6673934811591 17.2316886011198,53.6613940146887 17.2185716417436,53.6424681290096 17.2188627725109,53.5987859585823 17.221570996105,53.557344373748 17.2180300745752,53.5447132433727 17.2190256413875,53.4899248996613 17.2140640098801,53.4133356390444 17.2191757117935,53.3745260445819 17.2154242283351,53.3555221635339 17.2199285567752,53.3407627049203 17.2329916318333,53.337335979827 17.2468662055182,53.3414617118442 17.2614843988831,53.3464939694612 17.2688042007644,53.3680954988911 17.2862070609766,53.3708914925266 17.3044368875603,53.3624074228069 17.3188261770836,53.3408457299294 17.3244926117212,53.3127394005391 17.313786146466,53.2984191223436 17.2994913896907,53.2819112423453 17.274932108825,53.2675822623849 17.2661831105396,53.2405985698011 17.2596202845928,53.2292522489713 17.2594074161648,53.2184375366874 17.2640510229503,53.2063649533133 17.2778942718223,53.2059146222433 17.2904733095492,53.2193630663332 17.3113276673099,53.2394022643881 17.3287895552054,53.2815193150336 17.3529607395593,53.2938060606769 17.3626262675592,53.3110833691642 17.3647799505993,53.3147141446429 17.3682020232057,53.3155784609245 17.3829575262929,53.323321433409 17.3934881805661,53.3196250222885 17.4077232793871,53.306726428933 17.4214210060459,53.2838528144845 17.4288722751175,53.2574763253113 17.4223188986933,53.2429900362876 17.420834214738,53.2342443948302 17.4164277223108,53.2273317908702 17.4086275548016,53.2565313718648 17.3658641644997,52.9745924827323 17.2525853197983,52.984843095415 17.2193479123482,52.999074496676 17.1962335099226,53.0205831337837 17.1828606718376,53.043100939669 17.1806043563941,53.0575714515191 17.175188167068,53.0763327439646 17.1734543289349,53.0853267482288 17.1751204151322,53.0946138491382 17.1674232965725,53.1010574209602 17.1442739914299,53.1165477449184 17.124699846487,53.1300633487249 17.1194090335353,53.1510432305561 17.1223162281547,53.1600213763604 17.1203385364834,53.1660985384993 17.1145455017203,53.1795175759783 17.1139043140689,53.1839116355479 17.1084368817402,53.1826454679482 17.0792285036201,53.1917632611792 17.0702687142757,53.1978939738508 17.080052477889,53.2103622673934 17.0802861662393,53.2176470902304 17.0883006386535,53.2263363555172 17.0913276566611,53.2309507161942 17.0840723998219,53.2272443918922 17.0739763719769,53.2353291116219 17.0700084981895,53.2450736402505 17.0760981770581,53.2547937632091 17.0741294093557,53.2686730685468 17.0606508409238,53.3863486983556 17.0921163294725,53.3987223837785 17.0852185775127,53.4043229838116 17.0882046656859,53.4086168768171 17.09852848514,53.4223692432505 17.0977673942284,53.4475535129536 17.1001702107989,53.4561024415356 17.0983609212707,53.4674927155617 17.0899194586136,53.4812088221007 17.0966388418502,53.5117323727005 17.0957605466219,53.5210391787585 17.0925045075454,53.5352838988151 17.0962152912083,53.5351339788958 17.0845453992073,53.5405508885394 17.0720358365901,53.5539966727127 17.0659061858331,53.5560626828722 17.0575223938428,53.5753665704764 17.0424835473781,53.5890691419138 17.0400820222974,53.596179727064 17.028716634879,53.6061117861869 17.0240966307484,53.6191106313397 17.0039700792525,53.6219755591281 16.9926511353509,53.6284339281638 16.9900028985101,53.6355512537697 16.9796103774612,53.6387264587191 16.9521723283728,53.6295993859583 16.9397038589341,53.6370160895435 16.9338178941847,53.6333551415038 16.919353394597,53.6346753997748 16.9041912945753,53.6438515273 16.8995760556567,53.6582876045839 16.8968268642282,53.6633331670425 16.9016043146425,53.6761963476368 16.8924359745873,53.6564796959297 16.8704131799345,53.6708331838852 16.8609013392954,53.6734383125188 16.8492661950838,53.683248121309 16.8562472728582,53.6952491214712 16.858683228321,53.7109406835001 16.8568898738238,53.7165402858676 16.8661705217009,53.7262980225754 16.8686309072435,53.754728287116 16.8702802043016,53.7744445690117 16.8793481066439,53.8245692649732 16.8875929268594,53.8345569682934 16.8850863262514,53.859801478781 16.8903349513252,53.8684865529026 16.8946425333519,53.8910269760559 16.8968395336575,53.8994184910572 16.8938601433881,53.9190583431729 16.8996648483601,53.9331200334738 16.8975997375634,53.946359811689 16.898653438263,53.9488919313727 16.9097763903262,53.9615081245955 16.9121512319152,53.9644065567204 16.9085001094981,53.9757126361453 16.9135385051805,53.9790896632493 16.9224428047567,53.9907701543227 16.9286139591618,54.0050006206948 16.9291722684855,54.0115572358846 16.9397793797358,53.9991111224282 16.942271032655,53.9965168167289 16.9542108564961,53.9984212661602 16.9619312323732,54.009360713327 16.9745228485806,54.0275555288627 16.9850084098393,54.0484830069183 16.990828950095,54.0990072616984 16.9982601734863,54.146255147118 17.0063664024685,54.1884013904503 17.0127344278805,54.2179491293693 17.0162545798655,54.288696575478 17.0274982679906,54.341918296573 17.0316897681505,54.3394810429385 17.0532865288308,54.3420296783292 17.0611297539931,54.3316265609454 17.0642248219803,54.3205983168218 17.0620596955423,54.2986087029291 17.0531505822188,54.2749356449547 17.0543152171232,54.2681718308247 17.0506532870678,54.2491898469013 17.0532716302036,54.2387275312855 17.0717610220964,54.2335184422624 17.090759979966,54.2432687084464 17.098111528152,54.2544756250448 17.1009867482311,54.2573261263924 17.1075889511152,54.2651791601233 17.1115737047415,54.269797372398 17.1223002168863,54.2678642142944 17.1311820699552,54.2754722424394 17.1397571703852,54.3051923093605 17.1816712793552,54.2956604217455 17.2020846990975,54.281410374647 17.2045554003689,54.2796950193499 17.2126769404264,54.2941323834261 17.2249116276991,54.2962410048205 17.2490115069487,54.3075570833379 17.246014250337,54.3161534078258 17.2319024834728,54.3209066202708 17.2327582820497,54.3228112012221 17.2487549340234,54.3149205979886 17.2657249271423,54.2989925146391 17.2604674106444,54.2890175489326 17.2616256020981,54.2853202980322 17.2683059316176,54.2904173529812 17.2770173923312,54.2891411883231 17.2894447492353,54.2854421061579 17.2952907445055,54.2897385130626 17.3042646999342,54.2849693200102 17.3165830499782,54.3049482995579 17.3250383638969,54.3049921496272 17.3370022500973,54.3101471152306 17.3431582368418,54.3208991169093 17.3401543011274,54.3306068324161 17.348889417749,54.328029899255 17.3608184555843,54.3498397339335 17.3640473673101,54.3547346923736 17.3580254547748,54.3538137863553 17.3460495929237,54.3710128745194 17.335362096216,54.3841703201751 17.3321762578768,54.3932619605621 17.3228496310698,54.4121165409057 17.3184764925348,54.41683514964 17.3248343696144,54.4179288791555 17.3403809539426,54.4291013225838 17.3541683256386,54.4384980886349 17.3542889647882,54.4461936134858 17.3667716361368,54.4547082668546 17.3675100181084,54.461942388498 17.3626486907152,54.4741304887787 17.369855598914,54.4951119513884 17.370119834386,54.512116323299 17.3850811323603,54.5247739590573 17.3801172376013,54.5442848726058 17.381149654981,54.5536707810618 17.3860486769937,54.5793335056818 17.3829066438558,54.5966548171411 17.3976313736803,54.6286940745658 17.4056757738546,54.639292977886 17.4029031289065,54.6305834086636 17.4266339827413,54.6254933861438 17.4458210235288,54.6258353976599 17.4584314192187,54.6193204068271 17.4631115048723,54.6193088951347 17.4703984901142,54.6127862565292 17.4794511307398,54.6178304595637 17.4903825002186,54.6152720109076 17.5070237924173,54.6271740840006 17.5268656902998,54.6275164172852 17.5389972989193,54.6358229520044 17.5468602465519,54.6427009136416 17.5431315607886,54.6470575913315 17.532244669684,54.6636993198256 17.5290203946992,54.6705630002873 17.5350143676777))",Wilayat Salalah,ولاية صلالة
"POLYGON ((56.8848922287047 23.5964730407166,56.8777645206642 23.5978530453692,56.8579018197882 23.6188250942015,56.8697069163328 23.6428662224856,56.8630904783774 23.6529492883512,56.8523198295319 23.6513445898594,56.837708662909 23.6548097162609,56.8253490178493 23.628636281436,56.8066910324141 23.6222323803376,56.8111769123004 23.6455019401396,56.8084153466469 23.6810176083761,56.763387247019 23.6288327828902,56.667331457604 23.7069479633192,56.6495161053331 23.727741618394,56.5900527862972 23.7167430648257,56.5669245366057 23.6774027928617,56.5659146553283 23.6589533195302,56.5927062729867 23.6474799627038,56.599699150996 23.6236586706037,56.5807482466519 23.6144081701142,56.5890205236688 23.6023614101895,56.5693422813295 23.5884351864717,56.5769052839787 23.575272602902,56.5868366595159 23.5756656117063,56.6041445054678 23.5582641288564,56.5829814820682 23.5354524437455,56.5821823497219 23.5026692395139,56.5568653044212 23.4862639990812,56.5864089702656 23.4502206615106,56.5786542827293 23.4326171454959,56.5824543749168 23.4161975132628,56.5734298584468 23.4057963843117,56.5806829372253 23.3836212365197,56.5606982588578 23.3835663763382,56.551349879102 23.3777749651719,56.5576416640074 23.3636689257919,56.5504869848093 23.355865940678,56.4835895012901 23.3784306596902,56.4692526684279 23.3717531193742,56.4539275287672 23.3780416738995,56.4192742947264 23.3847977879979,56.2631127896109 23.4741173021943,56.2083120155417 23.4872800509741,56.1790339050576 23.4847705687005,56.1485011860388 23.4939850819043,56.0109662657225 23.4792860447887,55.975781252303 23.4981388754436,55.8851843571015 23.5133628277196,55.7622905011625 23.4706455691061,55.7082570786448 23.469054521229,55.6904625084701 23.436051834815,55.6826707170731 23.4028437629805,55.658966595819 23.3622815312256,55.531116910258 23.3356795997118,55.4173184319815 23.3830987964139,55.4016698859183 23.3923056601828,55.3557059287526 23.3085561575773,55.3479975781963 23.2929717089437,55.2990788662599 23.2068992153342,55.2803798640295 23.1769593719425,55.2519983675766 23.1418823010338,55.2364778888115 23.1190386812084,55.2324677511282 23.1104139007644,55.2314392318864 23.0853154669298,55.2256320696987 23.0724063766783,55.2303443580178 23.0555782311719,55.2301228350048 23.0479133828723,55.2185020024511 23.0332915810374,55.2165759645986 23.0262425425451,55.2173589284537 23.0096796430059,55.220512364654 22.9945239181812,55.2172889319598 22.9861202792977,55.2200242282497 22.9783423452461,55.2175637678394 22.9605979039768,55.218769482924 22.9519978592317,55.213639489917 22.9355560641407,55.2176895557448 22.9003247766392,55.2232598758169 22.8928897618457,55.2257278687695 22.8753487865436,55.2232455160681 22.8592752339215,55.218216129489 22.8509916242091,55.2219360553232 22.8326763430865,55.2265718967782 22.8251193986812,55.2236687960741 22.8172639357855,55.2280875640623 22.7915340410318,55.2207192810961 22.7649111617458,55.2157550332768 22.7271332998736,55.2083333182755 22.7083333504779,55.6666666728654 22.0000000373484,55.4439124493263 21.3373088530363,56.577367899338 21.4908794452847,56.6022469409291 21.6490577474757,56.6225688238349 21.6585618785817,56.6339462979413 21.671662627813,56.6361031497859 21.6923125125637,56.6294400774455 21.7064052354445,56.6139764292313 21.7237927934693,56.6358696174051 21.8667179688806,56.6396260452118 21.8878865502237,56.6550283885938 21.9871662411465,56.6571939028692 22.0045856866514,56.6708371484791 22.0931856024429,56.7026659379106 22.2374319992063,56.7356105180489 22.2502220111905,56.762836778117 22.2940622063036,56.7739113587372 22.3118855840309,56.7744479601071 22.3534560655595,56.7862432386579 22.4027187697778,56.786940139017 22.4703368349447,56.7986486023276 22.4717073038441,56.7977129778548 22.4806327363134,56.7871135066467 22.487152246743,56.7872951725845 22.5047701604025,56.7648775493956 22.5406902607666,56.7597455616434 22.5852141336849,56.7786437565569 22.6251572444698,56.7822537152524 22.6369585451552,56.8376363063073 22.6870180692113,56.8890389962391 22.7185187189212,56.9457195290254 22.7292208449242,56.9850586887522 22.7324124953675,56.9961539857765 22.7595632269188,56.990301019235 22.7758529274121,56.9525515667859 22.8082388722136,56.9392312277962 22.8031788424478,56.9053017778457 22.8303121139811,56.8860982313042 22.859134377095,56.8977012127194 22.8771171252853,56.8888055479081 22.8851274348799,56.8884489487416 22.8906727468172,56.9077768586653 22.8927282047229,56.9177720985311 22.9082105308374,56.9389730117577 22.9295652498818,56.9348290737217 22.954366638528,56.9226550939765 22.962636479535,56.946484281847 23.0318274979794,56.931644107119 23.0400317235076,56.915082597034 23.0439311272938,56.9130726674589 23.0488374384913,56.9213929694591 23.062449641667,56.929415571604 23.0677135637285,56.9574901031644 23.1163023606107,56.9299717622437 23.1456307864969,56.9313781645423 23.16547803008,56.9572868956513 23.1559383052667,56.963560369944 23.1565015695223,56.9590998319249 23.1836492792936,57.0244831848497 23.2001290237258,57.0779359578782 23.2145284396679,57.0779605682882 23.2569024115974,57.1237558968639 23.2851661132575,57.1431457064386 23.2892888655115,57.1398326019131 23.3008695446255,57.1188660853235 23.3117556827149,57.0833631221438 23.3187908089929,57.0714485620544 23.3323487359329,57.0887326857516 23.3712242339003,57.0570409947282 23.4119548306984,57.0226635116953 23.4407785693073,57.0073974767621 23.4514719633033,57.0205122736929 23.4668760729069,57.0781111618808 23.4896179497523,57.0939741276902 23.5072933756842,57.0360308316768 23.547668422976,57.0041785903287 23.5635385770995,56.9866105451378 23.5412368579328,56.959710611883 23.5333182228394,56.9485447722418 23.5317235001861,56.9255450165945 23.5443881516878,56.9172358517373 23.5575858518087,56.9184561766945 23.5904156845971,56.8848922287047 23.5964730407166))",Wilayat Ibri,ولاية عبري
"POLYGON ((58.8860903179293 22.7798809746318,58.8730845940949 22.7932906772854,58.8706335185412 22.804187398114,58.8742916323772 22.8178049480439,58.8919602805574 22.8312000744698,58.8838302223511 22.8421868771717,58.8735971664229 22.8418764544795,58.8576323670289 22.8595890680017,58.8428701580077 22.8602890261172,58.8421195131631 22.8815302446034,58.8392093412024 22.8881876718722,58.8178715081212 22.9026763124739,58.8083995701631 22.9028250541882,58.7967811513867 22.9100819001681,58.7729697692738 22.9137472235735,58.756265039337 22.9121244708217,58.7377486835132 22.9152360173174,58.7233040179018 22.9085869322208,58.724694460394 22.9047841648132,58.718843406408 22.8897675770006,58.7036104929965 22.8579670015919,58.6669929057621 22.8465817145854,58.6585874777142 22.8419756288732,58.6497226088593 22.8442222660731,58.6395058226614 22.8332905539742,58.6255223069169 22.8324202724074,58.6131164650749 22.8213537507427,58.5828347399612 22.8104101387205,58.5797238897254 22.8000681518259,58.5719609689433 22.7883906639716,58.5721416671839 22.7761130922031,58.5754575075161 22.7704064748496,58.5756001355032 22.7557856389463,58.5730254416173 22.7369445713559,58.5741077488173 22.7253388506407,58.5830114168743 22.7197886134275,58.5809028182967 22.7097510450978,58.5865463686422 22.7070301173093,58.6082226606508 22.6670895181534,58.6202680824847 22.6515293299689,58.61480384898 22.6424329831683,58.6171386610115 22.6339316530866,58.5897173769806 22.5989381902599,58.5840400854526 22.5902870089286,58.5899867348593 22.5812796104578,58.6069879415709 22.5684764401063,58.6094632432081 22.5588405845308,58.6002239133616 22.5568303878871,58.5927083792676 22.564113376626,58.5681486434628 22.5704276958206,58.5560364801998 22.5783806425982,58.4894146577752 22.5701623042403,58.4661677184414 22.5657174338085,58.4530163897223 22.5661043858932,58.4338168206208 22.5746634185479,58.4210431379664 22.5700577617672,58.4276236205336 22.5561710554946,58.4376725421565 22.5457037882681,58.4579144084094 22.5389176093836,58.4652639666239 22.5212609378503,58.4800907911352 22.4792831667778,58.4977881980113 22.4637133814487,58.5079099000624 22.4473161041588,58.5004256404748 22.4096943718055,58.4618485436933 22.3817788714014,58.4502183185346 22.3616858862897,58.4363115682587 22.353236494051,58.4342420881067 22.3399460162336,58.4449819339684 22.3278429074518,58.4731424346003 22.3231298443261,58.5032405217862 22.3122978730999,58.5044859247937 22.2892430839158,58.5136341545529 22.2652847912012,58.5181552632715 22.2352683770526,58.5123469298374 22.1984513556061,58.5022879082749 22.1632646297161,58.5030827707285 22.1455413559629,58.5330496789184 22.1333534559499,58.5598551466618 22.2083222242976,58.5985583475404 22.2377579593309,58.6082775207804 22.2754379613968,58.6162724250798 22.3115412117055,58.6189698412689 22.3333603283569,58.6331863762336 22.3440142412413,58.654326646928 22.3441835344403,58.6546990612202 22.3668261622785,58.6743071448705 22.4108940598947,58.6948394725484 22.4417317825138,58.6998936431196 22.4604269831594,58.7026473422057 22.4800672826316,58.7132791891619 22.4970831688583,58.7425552697682 22.5221941696615,58.7377472635547 22.5390369182285,58.7319951077148 22.5511203371592,58.7403850564879 22.5683235812447,58.7462349934191 22.5738548254213,58.7443047185737 22.5830532741107,58.7409073131827 22.6235643621208,58.745467864295 22.640068108653,58.7558822885958 22.6516967244106,58.7839180006403 22.6758382121223,58.7958228357578 22.6784590995581,58.8118352639593 22.6774524835235,58.8269206925061 22.6737009092377,58.841729599172 22.6747802402113,58.8619795249534 22.6823419822836,58.8917219938934 22.7032409712322,58.9291735128941 22.7053678973458,58.9346368834124 22.7118203971132,58.9364193046775 22.7210013925068,58.9058120061774 22.739391154484,58.8865129510536 22.7589204008722,58.8860903179293 22.7798809746318))",Wilayat Al Qabil,ولاية القابل
"POLYGON ((58.0687978254054 23.7135745793987,58.0458281124629 23.7144723994631,58.0170032696487 23.7135802004985,57.9559000593766 23.7082184225839,57.9260776556469 23.7080103647876,57.8865072523543 23.7109353384698,57.8566668307246 23.7201899364078,57.8213702098385 23.7399009683482,57.8056302019496 23.751669203884,57.7927725082996 23.7686794352536,57.7911104805638 23.7823984378588,57.7701962990879 23.7730807264905,57.7452828285943 23.7682027390839,57.7183784849034 23.7693102827304,57.7206573329982 23.7579930953636,57.7177334501611 23.7459156072721,57.7100203336916 23.7409557404613,57.7062917204027 23.7291241626379,57.7097746540638 23.7227570626611,57.706691809966 23.7069414694753,57.7015909648506 23.6936203977761,57.6901425416215 23.6508111866167,57.6626335609093 23.609683169844,57.6455202257619 23.5354355570249,57.6904054401984 23.5383397873566,57.7163510517146 23.5869053670187,57.7346941486798 23.5919576099111,57.8517497080017 23.5757797684817,57.880732222366 23.5595300568129,57.9923532749528 23.5821922588092,58.0085388161426 23.5919040394889,58.0278021330441 23.5926053969556,58.0535001300214 23.5821584504815,58.0816830738052 23.5628765732803,58.0954386276463 23.5803891506245,58.0924556065835 23.6047573186043,58.0870370644335 23.6097311157798,58.0865196381516 23.6198687472315,58.0897699333467 23.6319932695804,58.0753441027865 23.6513799411948,58.0741977322513 23.6570822656575,58.0864536473341 23.6687285490993,58.0778072695916 23.677126253309,58.0782011980285 23.690869463789,58.0645524901368 23.6932460825867,58.064149894467 23.7005440872851,58.0687978254054 23.7135745793987))",Wilayat Barka,ولاية بركاء
"POLYGON ((58.041880705831 21.3517685337677,58.0183138339252 21.4746774863853,58.0145450389967 21.4975344819953,58.0140813948249 21.5176959602389,58.0812254167827 21.5850850122039,58.0512449770805 21.6305955535301,58.0292212497345 21.6612086922124,58.015357510206 21.7002713751336,57.9439209464011 21.7003445062584,57.9392798354492 21.7240566881746,57.9675182052809 21.7373212319654,57.9670375247868 21.7724415710174,57.9437345283352 21.8285313108614,57.9197632173897 21.8589746799383,57.8823735434358 21.9079636277549,57.8618258011444 21.9581477256949,57.8399912112635 22.00544379027,57.8317801078301 22.0258741714211,57.8158351688434 22.0438331587693,57.7865405917639 22.0727502739145,57.7636217748654 22.0925755597166,57.7321485565712 22.0922716470253,57.7273646796641 22.0817729909505,57.6679691275807 22.0640553341978,57.6623544587289 22.0878520076207,57.6940299900165 22.1089189323367,57.7122354734107 22.113348083222,57.7115601985547 22.143694602983,57.7079918786056 22.1565414688159,57.7122144883978 22.1681812631098,57.7176454486866 22.2093141989613,57.8274075347575 22.3257127414043,57.9061786237177 22.4102653608332,57.9045408426286 22.4878387001794,57.8785060531634 22.4855646761178,57.8675006468121 22.4865379287457,57.8549500761089 22.4920868979524,57.8560468289483 22.5105368209029,57.8625786484723 22.5172629688844,57.8939798742437 22.5373745276702,57.9041180311541 22.5476842769221,57.90430268359 22.603321718951,57.6744523732107 22.5137949020557,57.6759015291704 22.4996876378843,57.7020623407205 22.4721822026744,57.7005195628586 22.4605613950939,57.6862719150105 22.4521483058827,57.6512890758618 22.452293269284,57.6377532544282 22.4596392336495,57.6306030942587 22.4726745201264,57.632788068992 22.4868555899997,57.6263304123396 22.4949944380171,57.6365977437997 22.5347363600622,57.6290960608466 22.5949951799129,57.5597431958942 22.5437727907137,57.5283106520874 22.5667773497906,57.5260935933885 22.5814276801781,57.5110075378977 22.584367006355,57.5130171774783 22.5779652502905,57.3832967815503 22.5502026199542,57.3875149441882 22.5594459308724,57.3800724845484 22.5631553882492,57.3648990594252 22.5558071468251,57.3420319232345 22.5505505785692,57.3305893732544 22.543883273411,57.3303610021942 22.5388399480485,57.3167473924131 22.5359146574757,57.2405508589168 22.4884784600897,57.2107083976502 22.4604932020885,57.1878978133028 22.4567076816885,57.1325869331343 22.4892925121657,57.1013375710192 22.4604857861491,57.080678491111 22.3440863340711,57.0174573355013 22.3061653155684,57.0045990750416 22.2921832595225,57.0038661237096 22.2665827974693,56.9986535579405 22.2411066630328,56.9842370853745 22.2412150931346,56.9515337082296 22.2472972381213,56.9182809820048 22.2559094318221,56.762836778117 22.2940622063036,56.7356105180489 22.2502220111905,56.7026659379106 22.2374319992063,56.6708371484791 22.0931856024429,56.6571939028692 22.0045856866514,56.6550283885938 21.9871662411465,56.6396260452118 21.8878865502237,56.6358696174051 21.8667179688806,56.6139764292313 21.7237927934693,56.6294400774455 21.7064052354445,56.6361031497859 21.6923125125637,56.6339462979413 21.671662627813,56.6225688238349 21.6585618785817,56.6022469409291 21.6490577474757,56.577367899338 21.4908794452847,56.5262051183743 21.3277858407854,56.6288489946401 21.2730143513206,56.6315664404592 21.2655798309765,56.6518802274495 21.2298853091513,56.6861257076206 21.2212003416346,56.7075739395412 21.2359829222017,57.1221718176992 21.0599769344571,57.3391767426874 21.0115322059444,57.4665875616156 20.989135143368,57.9851096563674 20.8977971391021,57.9946014243532 20.9407148689552,57.9910575043536 21.0496791161221,58.0140287042868 21.1143229631068,58.0387860776851 21.1401323409548,58.070465914996 21.2024710729628,58.041880705831 21.3517685337677))",Wilayat Adam,ولاية أدم
"POLYGON ((56.4865396656246 19.0938157204497,56.4705965934749 19.0950268283152,56.455891366393 19.090465138602,56.4393388448401 19.0992274675466,56.4282124695064 19.1010317462257,56.4122801833183 19.0945469181164,56.4002399026315 19.0816387684353,56.3015591597526 18.9793905976889,56.3000658008617 18.9785705896532,56.2475812029582 18.9853836513755,56.1940951797382 19.0379639728825,56.159302034385 19.0947780549616,56.1572334900845 19.1053461727701,56.1469182002006 19.1178751056816,56.1095068726772 19.1172814538915,56.0916147462422 19.0883767890257,56.1015368152674 19.0551682353469,56.0852670095965 19.0044544104995,56.0784617047 18.9724367643168,56.079446577496 18.9578113732898,56.0777085363308 18.9448936318646,56.0978320989593 18.9028226016464,56.1269270736877 18.8719792241844,56.1273847805011 18.7833368111428,56.0789019530524 18.7857850809901,56.0509643973851 18.7910061213276,56.0180136869433 18.7992392998394,56.004876752186 18.7991482680057,55.9655442654266 18.7877119814003,55.9186973266928 18.7566464331016,55.8402280132996 18.7163673047502,55.8565817421901 18.6911301010414,55.7663842739647 18.5989966326859,55.8413951844763 18.4897889958427,55.8515155336813 18.4920628717873,55.868387156205 18.4903662564688,55.8828463880479 18.4969635441073,55.9270805938945 18.5090223145744,55.9684209435662 18.5182865053955,55.9858954350691 18.5152453306629,55.9979481760327 18.5073924624753,56.0003783363524 18.4841592644063,55.9946283204056 18.4777204910562,55.9694533515313 18.4725950319863,55.958120296298 18.4738509281263,55.9445406989223 18.4698909425214,55.946630604823 18.4528472131174,55.951247638415 18.4446293580058,55.9670214285953 18.4419598478503,56.0149679382374 18.4462205857403,56.0237167595048 18.4326668676184,56.3450819376393 17.9329781413001,56.3536691272746 17.9210449091626,56.3555743606668 17.9312754903583,56.3503076435691 17.9425478324122,56.3537631572138 17.9579604778982,56.3615164115525 17.9676152199254,56.3731815309637 17.975482609932,56.3864963488758 17.9802928456185,56.3941152113598 17.9889652645461,56.4069821848551 17.9960447180096,56.4138441364719 18.0039876238001,56.4274193583628 18.0144674159402,56.4312607787281 18.0211207291812,56.429633776566 18.0388309066236,56.43687264126 18.0516321933399,56.4479444548776 18.0611429936759,56.4837656822037 18.0830174910906,56.5058586124204 18.0918401967245,56.5110132324664 18.0955409511909,56.5190361872514 18.1088312325606,56.5289876719607 18.1173836096021,56.5445132138655 18.121889921371,56.5509731536036 18.126664834811,56.5485860869483 18.1584453455399,56.5441805616074 18.1669076302169,56.5441903988401 18.1785703006008,56.5490531907369 18.1853775392968,56.5580154834384 18.2267066942277,56.5865534989496 18.2710114439862,56.5903469794251 18.2849241407857,56.5994289125197 18.2996810912709,56.6037821811644 18.3260262720271,56.6082587804031 18.340719129821,56.6064367034723 18.3605224574506,56.6091687988327 18.3964159569927,56.6231749020338 18.4274323279552,56.6332610428495 18.4455089828535,56.634115675165 18.4539380883062,56.6312698144998 18.4720972557283,56.6262631899218 18.5296309061792,56.6327749574241 18.5477910359949,56.6294390982437 18.5536101103416,56.6361289907321 18.5747814189934,56.6583373756367 18.5982130154565,56.6692125945378 18.6061611547999,56.6859276221376 18.6247669404273,56.6959990348066 18.6388882849235,56.7213489418045 18.6679811307222,56.7393857038405 18.6861174159625,56.7304865372792 18.6948352731705,56.7258162668408 18.7073344536025,56.7279049354262 18.7336168010872,56.7027759237275 18.7579149129255,56.6920403287071 18.7704646208975,56.6886954373369 18.7856538729299,56.6831526076104 18.7982161021059,56.6711630370842 18.8120717143793,56.6582339708292 18.8198966243302,56.6443525575591 18.8243127110341,56.6329680366341 18.8245425769934,56.6183372888415 18.8289552317193,56.6143259136655 18.8349694649941,56.6102024668205 18.8535604132547,56.5987511151757 18.8758583969501,56.5962761385984 18.8977605347645,56.5953756307144 19.0277431016628,56.5820610094222 19.0623765655521,56.4944825157537 19.0906541909349,56.4865396656246 19.0938157204497))",Wilayat Al Jazir,ولاية الجازر
"POLYGON ((56.5611249232296 24.5790028568444,56.54092231362 24.6098447674026,56.5260295545943 24.6390240254726,56.5080118452982 24.6685918025631,56.4958903891281 24.6930231336764,56.4908434670345 24.6996364311049,56.4762351206721 24.7319575432525,56.4678621287784 24.762976176063,56.4546273459447 24.7988750975724,56.4394187406282 24.8259781766062,56.4268302807902 24.8421826559235,56.4153060532109 24.8711917383739,56.4113735003761 24.8750732952359,56.4035420914516 24.8988353083585,56.3926045725462 24.9214968142535,56.3831984916728 24.9490822649038,56.3747107331521 24.980440067927,56.3512321319085 24.9762371123552,56.3433904863637 24.9718206542258,56.3235783974135 24.9723381006897,56.3412027924687 24.9420563603122,56.3500661194798 24.9339514058124,56.3389151034108 24.9143848318458,56.3260902321324 24.8981713272159,56.3053686464714 24.8842196269019,56.2805960556567 24.8842133649081,56.2806535673269 24.8750340402437,56.2591324368139 24.8599502879646,56.2058829762108 24.8502575673982,56.2012181333435 24.7843983083917,56.1893392386152 24.7781721670329,56.1902334889336 24.7699433578057,56.2017592239465 24.7601491945028,56.2012875692826 24.749551547286,56.2176880454103 24.7359629126459,56.2105150950118 24.7189235416316,56.20776927219 24.7054801526812,56.202286165506 24.6986750552714,56.2076150307853 24.6872456037495,56.1982916298347 24.6699479900005,56.2064895005422 24.6521272499988,56.2034970164724 24.6353560295668,56.2365390531043 24.6301300041053,56.2484956915338 24.6052082845602,56.2333464734511 24.5988863904977,56.2097985052325 24.6102247401222,56.1842378596012 24.6138157580224,56.1833670737494 24.6027228200743,56.1760236131247 24.5929498581652,56.1756850005439 24.5829685980281,56.1887000550963 24.5484193102135,56.1837813647145 24.5387829229006,56.1940279816967 24.5362507248792,56.2376160493442 24.5408889023225,56.2753173397952 24.5464142738584,56.3135837026625 24.5498057807124,56.3669107691476 24.539814788067,56.3716645984331 24.5737554743686,56.3712525263257 24.5904284294458,56.3884509719013 24.6043321762625,56.4059805354049 24.6011696791035,56.4124642413297 24.5949702991384,56.4546593496852 24.5630348716339,56.471676335606 24.5529461969283,56.5105302293228 24.5508219456116,56.5408350192318 24.563046489019,56.5515917471391 24.5801493215928,56.5611249232296 24.5790028568444))",Wilayat Shinas,ولاية شناص
"POLYGON ((59.8232483508265 22.360452949277,59.7916656907279 22.3605174280422,59.7135054691501 22.3553767751266,59.704631130374 22.3677845673031,59.6942466208153 22.3646565192907,59.6985990644119 22.3506996834679,59.7088911805478 22.3310394039781,59.7122808726534 22.3076848201277,59.6605145307538 22.2780438503401,59.6378774948486 22.2733074820527,59.6151298746662 22.2732768004873,59.5777099755223 22.2471363312277,59.5522234586209 22.2419328688639,59.5486036853776 22.2366888872238,59.5519151226396 22.2204718358326,59.5441351084601 22.2136679050294,59.5284380625384 22.2077387552054,59.4921926447481 22.2065160691032,59.4755842401944 22.2074151487596,59.4740102905363 22.2006633615444,59.4846353173464 22.1762019551284,59.4676571066379 22.1517449089695,59.4261958319379 22.1251826007808,59.4118880387445 22.1176576532123,59.4108535489606 22.1032816316995,59.4127104564645 22.0701978838535,59.3998872173722 22.0657807106554,59.3567964875126 22.0606486671379,59.3308747201718 22.0638809875231,59.324208954164 22.0578949048719,59.3165102584095 22.0571265182572,59.3042320411142 22.0434290087628,59.2916280114146 22.0428368958798,59.2851588405814 22.0382162913686,59.2847505185452 22.0267642274793,59.277803641555 22.0254535814637,59.2616549564621 22.014719391487,59.2484297430508 21.9967989545244,59.228471805024 21.9980175688069,59.2100409540596 21.986664211126,59.2117559482254 21.9692407970845,59.2098146714891 21.9521543351106,59.2175499186554 21.9476816164137,59.2310524004413 21.9527408475912,59.2570779326353 21.9698585896596,59.2669152463076 21.970014212681,59.2719545044043 21.9629552142052,59.2569188722626 21.9499119638339,59.254398953735 21.9332015336058,59.2558435735687 21.907324952379,59.2823257995707 21.8536224208283,59.2876678392423 21.7990484649778,59.2870791773548 21.7619519081237,59.2704572264111 21.6766813186801,59.263633112307 21.6676656282726,59.2494830933009 21.6612910939552,59.2125107234575 21.66651304944,59.1752751205448 21.6544082680953,59.1749684921411 21.6339453665669,59.1931691790532 21.6010088580843,59.2250956539978 21.5806406246003,59.2383411352088 21.5750075511621,59.2473636107754 21.5764666208211,59.2576432383956 21.572961167066,59.2751298305098 21.5456424560951,59.272307009337 21.505121193385,59.2571968518052 21.4769991642926,59.2577805667232 21.4743387452659,59.2445986161832 21.4535418106454,59.2403359439641 21.4426818720213,59.2052519175106 21.415781910439,59.0849490585331 21.3438158781291,59.0377677446359 21.3349484581808,58.9990780844017 21.3322636102079,58.9786721550959 21.3322057235353,58.9708013461071 21.3231995073333,58.9688792567802 21.3148045828243,58.9763343375928 21.2987081929137,59.0336917217238 21.2830373958973,59.0199964638301 21.2643067708461,58.9876202022621 21.2300498668939,58.9113066781793 21.1726683136766,58.8203522081033 21.1484771149746,58.7726505963806 21.0783795826631,58.7366961758017 20.9716858835556,58.7967450851588 20.9709184766572,58.7968835240989 20.9797137075127,58.8014997732341 20.9918764552071,58.8149440907022 21.0093036613535,58.8377470871983 21.0419754125787,58.8315697311502 21.047196261012,58.8555298407118 21.0811655141048,58.8642511792479 21.0768367784424,58.898842353074 21.1138848381537,58.9214471207734 21.1393135656302,58.9310897325139 21.1479452798178,58.9359476114182 21.1632601635444,58.9435489146352 21.166446597102,58.9450879610454 21.156961044257,58.9683304912961 21.1765279721381,58.9741856685618 21.1850747974604,58.9956136769845 21.209338734285,58.9999887867596 21.2163652657028,59.0156552093212 21.2316408356765,59.0123595036668 21.2391093327021,59.029203241875 21.2454714187237,59.057535784808 21.2690801854635,59.112348342781 21.3091017444302,59.1042333005722 21.3138118499852,59.1048265563451 21.3244861476205,59.1134695894126 21.3191322234391,59.1266189516903 21.319634815019,59.1457457033332 21.3316305140923,59.1498182897531 21.3364075626981,59.1863377837123 21.3652898857173,59.197386827063 21.3708040734112,59.2708408343722 21.3972668446253,59.2994928296102 21.4097211776973,59.2982748941308 21.4140775158998,59.3064748045946 21.4263543815851,59.2891049285536 21.4233147156109,59.2847994904197 21.4276632647131,59.2895670993758 21.4395898689554,59.2893576224467 21.4528518816565,59.2988522942195 21.4606185922988,59.3054853765054 21.4453183818332,59.3126627505911 21.4352266158384,59.3335177082995 21.435379622278,59.3406392615121 21.4412027631222,59.3419779240712 21.4569056608148,59.3434962699273 21.4653752926212,59.3499088866393 21.4750818716371,59.3830214198801 21.5128297497946,59.3794864779717 21.5159325775689,59.3828665735112 21.5285486231403,59.3983074574739 21.5465590648775,59.4192500092317 21.5783611511334,59.4282638567566 21.598256363551,59.4400774818911 21.6118165753498,59.4600544599042 21.6431728795703,59.4563408031071 21.6564267128592,59.4664200474546 21.6762980726178,59.4795527664933 21.6925138477059,59.4858810768417 21.7049937518901,59.48762294954 21.7167793505593,59.4833063530619 21.7254100949168,59.4857795529032 21.7387052243351,59.4922556490672 21.7549509389271,59.4981082596464 21.7637783396997,59.5175070586176 21.7857501297878,59.5568539382315 21.8251088112631,59.57571633588 21.8401936844576,59.571303593905 21.8513431255676,59.5764323404022 21.8683119466422,59.6075187887088 21.9063030483707,59.6453785756461 21.9353116071203,59.6528351471957 21.9485689690936,59.6452000219929 21.9613508471859,59.6464619330089 21.9706459681753,59.6576983821505 21.9895339539424,59.6593626509036 22.0003753051232,59.6684421388648 22.0153705216319,59.6746900971624 22.0368210950664,59.6696009451095 22.0442296371334,59.6749485411885 22.0662865099104,59.6912970362955 22.088955319841,59.7041541641701 22.0991355726035,59.7128589861262 22.1146207633358,59.7271622094151 22.1307032800797,59.7396788765037 22.1513961044454,59.7634327702686 22.1729178502542,59.7672859293656 22.1866233314512,59.7733873752125 22.198506649634,59.7970384660572 22.2186825578167,59.8097242029619 22.2260358286774,59.8071330945251 22.232448716585,59.8103889199523 22.2424082526972,59.8106858208108 22.2558928421742,59.8173805083865 22.2779133504907,59.823583231767 22.2919385049523,59.8213199830985 22.3178167178643,59.8227651709921 22.3237060705755,59.8154807802549 22.336799251108,59.8232483508265 22.360452949277),(59.7133277186826 22.2779290011056,59.7224363943284 22.2768438444484,59.7288471992103 22.251564918983,59.7358872356286 22.2442447961554,59.733743193385 22.2390286729475,59.7159290028346 22.2383312845649,59.7055466821681 22.2346105308068,59.7037200790295 22.2407988114637,59.6932525817998 22.2502908738251,59.6867521258682 22.243186204368,59.6816733800669 22.2473544630944,59.6756702559208 22.2622570500416,59.690184334102 22.2645247250681,59.6955544648458 22.2705691655549,59.7133277186826 22.2779290011056))",Wilayat Jaalan Bani Bu Ali,ولاية جعلان بني بو علي
"POLYGON ((58.2450239112885 23.4543713335279,58.2311261335369 23.4590350237451,58.2303666073906 23.463611508124,58.1881570766493 23.4748219797359,58.1835042052094 23.4733763968563,58.1632584525037 23.4784061494495,58.1497816159235 23.4946910270113,58.0766447333544 23.5007623240994,58.0609281457484 23.51297899983,58.0609506795656 23.4743454336585,58.0431701843931 23.4338248491112,58.0740104403202 23.3891355451027,58.0773081063557 23.3606179020888,58.1004858123198 23.364324459516,58.107161552849 23.3785767524944,58.1123327711566 23.3733224629356,58.1263357888263 23.3766047862114,58.1305474514014 23.3687317329282,58.1544214135403 23.3369209299095,58.1676475320334 23.3374564703384,58.2068285201202 23.3500324030617,58.2132660634493 23.3426308256966,58.2129665615083 23.3210629188753,58.1899157345405 23.2791089074749,58.2209137728906 23.2313950833118,58.2617015721919 23.2191237709741,58.2711291315975 23.1723047973153,58.2952992662861 23.1191718154691,58.2564145969243 23.0755949816373,58.2346219933729 23.0642630120859,58.2303411890025 23.0523692863411,58.2965205679133 23.062465423235,58.3134342280881 23.0916526960364,58.3469474898399 23.1010874746293,58.3587297362814 23.1058299505726,58.3892968043697 23.1129980902838,58.3902425127831 23.1232264317192,58.3758876507609 23.1289682572517,58.3706095727406 23.134726495066,58.3426395558817 23.1430943773073,58.3424045565356 23.1764488355156,58.3491418058643 23.2159816571924,58.38338684108 23.2164818301514,58.3675820218537 23.2285720096729,58.3573732076725 23.2482179489343,58.374533190659 23.2514838282314,58.3609041939617 23.2660065714797,58.340132360524 23.2711528432161,58.3297494310354 23.3078768010933,58.3374742039902 23.3168859046639,58.3038883830302 23.3431774662158,58.3103629333383 23.3689490051002,58.3065872602882 23.3785487103259,58.2826059172647 23.4007841401843,58.2669696902108 23.4189257150644,58.251585954932 23.4271185147935,58.2450239112885 23.4543713335279))",Wilayat Bidbid,ولاية بدبد
"POLYGON ((57.058891250751 24.0224231987734,57.0336946356391 24.0437381773995,57.0227505774827 24.0489233932247,57.0016286624111 24.0636036564801,56.9554898033645 24.1004881040173,56.9321281869451 24.1230264749354,56.903152881623 24.1561290824455,56.8904713942518 24.173782575876,56.8727692626823 24.202383281479,56.862285281371 24.2126079797327,56.8414913653767 24.2393476107999,56.8302897859773 24.2283450130693,56.816861202911 24.2313942084522,56.8093952838272 24.2238310256967,56.7864522319653 24.210763587348,56.6693598797609 24.1790418303609,56.6036011852927 24.0940778989977,56.592306437568 24.0540718132166,56.5864121953945 24.0385411519884,56.5717893424014 24.0392790543121,56.5596722686423 24.0105396001834,56.5556043910468 24.0077093546925,56.6093817907965 23.9872646680539,56.6559944887482 23.9359631618412,56.6651997178926 23.9622883901113,56.6910543491704 23.9839155317281,56.723218540988 23.9764822427098,56.7355672040349 23.9598981000461,56.7747578380811 23.9680022600898,56.7803443402806 23.9674135421636,56.8228981109326 23.922873171815,56.8045857476312 23.8747226205568,56.8260396159744 23.8450922992754,56.7772425792622 23.7905373796658,56.7358414397874 23.7768046582167,56.7291382683574 23.7785679591413,56.7226791319721 23.786683712279,56.7114142195637 23.7896935502149,56.6926186893222 23.7353882562129,56.6477307172913 23.7528183475121,56.6401329881716 23.769023072177,56.6539332483305 23.7875218495692,56.6321682161665 23.8031143046281,56.5701032325482 23.778289873231,56.5606638530844 23.7785523401547,56.5498596450383 23.7831032543773,56.5673795941769 23.7551589952148,56.5900527862972 23.7167430648257,56.6495161053331 23.727741618394,56.667331457604 23.7069479633192,56.763387247019 23.6288327828902,56.8084153466469 23.6810176083761,56.8111769123004 23.6455019401396,56.8066910324141 23.6222323803376,56.8253490178493 23.628636281436,56.837708662909 23.6548097162609,56.8523198295319 23.6513445898594,56.8630904783774 23.6529492883512,56.8697069163328 23.6428662224856,56.8579018197882 23.6188250942015,56.8777645206642 23.5978530453692,56.8848922287047 23.5964730407166,56.8927118544688 23.6163858174042,56.8901362341169 23.6839336254225,56.8993728424919 23.7137135523303,56.8998612324199 23.7232471551562,56.9077360266087 23.7666250903258,56.9153337080125 23.8016187266885,56.9485052787326 23.8728271202045,56.9381574569653 23.893084118321,56.8614418462245 23.8940758614896,56.8716274186591 23.9191181815662,56.8826860868881 23.9527476365771,56.8963226418863 23.9667527877276,56.8969042991333 23.9717925220927,56.9667911376202 24.0212096858126,56.9839253396404 24.0294505330206,56.9969828300034 24.0444363236558,57.020981315412 24.0337904790356,57.0462707406998 24.0121700110424,57.058891250751 24.0224231987734))",Wilayat Saham,ولاية صحم
"POLYGON ((56.4251519045391 25.9296128209767,56.4217143512012 25.9367509632418,56.4118504363211 25.9377984879004,56.4020221364435 25.9461760032619,56.3947859069078 25.9472857986561,56.3765818857828 25.9400710405254,56.3711245865737 25.9323467576518,56.3645616141125 25.9153620235197,56.3571379171061 25.9131041151726,56.3491028255415 25.917920976859,56.3359559583236 25.9139989377279,56.3349562960548 25.9030571080117,56.3261930340355 25.8916192868664,56.3160189954004 25.8839122131211,56.310777736977 25.8642006006702,56.2986293043029 25.8475115662234,56.2804926950215 25.8412040210082,56.2798420399877 25.8552601978985,56.2636878714708 25.8535643079505,56.2616285010419 25.8597061412811,56.2363265904557 25.8606865431743,56.2301632152982 25.8628697908512,56.2289421983578 25.8777155637139,56.2204107418475 25.8671836549533,56.2039551728054 25.8756452821828,56.1983194575243 25.8859230685461,56.192628234753 25.8910078991936,56.1784278933725 25.89317130609,56.1693357165655 25.8871871997524,56.1597756757912 25.8755113011379,56.1641913466512 25.8650084930438,56.1629637956467 25.8579223451405,56.152655537305 25.8480295008312,56.1509009036678 25.8408137631896,56.1415849493641 25.8278649731595,56.141405616227 25.8126131708173,56.1548814929511 25.7973420099602,56.1567341417554 25.7610360214828,56.1604321329719 25.7555674270737,56.167700064207 25.7256489901927,56.1586049218817 25.6893428595103,56.1774826635266 25.6177095220603,56.202969665597 25.6191510240563,56.2155490961691 25.6160586558016,56.2284166254713 25.6098785107365,56.253351321678 25.6022964855257,56.266361529461 25.6064528804109,56.2594260390768 25.6182827967135,56.2709358306857 25.6258949485712,56.2688185766517 25.6338708215807,56.2692122879486 25.6577809703205,56.272335588639 25.6729979715612,56.2827648340957 25.6815541977487,56.2783354131986 25.6909937309784,56.2818450430002 25.6988409683563,56.2739129645475 25.7025652102078,56.2759977061045 25.7140313756746,56.3002897635693 25.7434174089499,56.311451620148 25.75040591781,56.3209980548592 25.7451486400881,56.3292365393435 25.7500767129574,56.3481570832464 25.7793514248662,56.3510129050668 25.7889120005102,56.3591863591811 25.7960016572474,56.3605503189578 25.8030244156461,56.3705432610745 25.8077243052238,56.3672906895299 25.8170576033744,56.3727277865616 25.8286025796158,56.3617303217923 25.8349176615489,56.3824859170026 25.8385621932137,56.3848103317635 25.8455665184067,56.3725215135221 25.8517849130963,56.3769478531055 25.8613085253426,56.3891812980431 25.8572684249147,56.3992112644855 25.8678264054678,56.404475161644 25.8799326919771,56.4005345646211 25.8833728524837,56.4089499595876 25.8982327814042,56.3952240425748 25.9012652099147,56.392435585193 25.9219229449153,56.3959283598569 25.9354320723465,56.4035669137504 25.931645718667,56.4251519045391 25.9296128209767))",Wilayat Daba,ولاية دبا
"POLYGON ((58.841729599172 22.6747802402113,58.8269206925061 22.6737009092377,58.8118352639593 22.6774524835235,58.7958228357578 22.6784590995581,58.7839180006403 22.6758382121223,58.7558822885958 22.6516967244106,58.745467864295 22.640068108653,58.7409073131827 22.6235643621208,58.7443047185737 22.5830532741107,58.7462349934191 22.5738548254213,58.7403850564879 22.5683235812447,58.7319951077148 22.5511203371592,58.7377472635547 22.5390369182285,58.7425552697682 22.5221941696615,58.7132791891619 22.4970831688583,58.7026473422057 22.4800672826316,58.6998936431196 22.4604269831594,58.6948394725484 22.4417317825138,58.6743071448705 22.4108940598947,58.6546990612202 22.3668261622785,58.654326646928 22.3441835344403,58.6331863762336 22.3440142412413,58.6189698412689 22.3333603283569,58.6162724250798 22.3115412117055,58.6082775207804 22.2754379613968,58.5985583475404 22.2377579593309,58.5598551466618 22.2083222242976,58.5330496789184 22.1333534559499,58.6253710632449 22.1002084916842,58.627162210127 22.0685033509303,58.6349931469328 22.0125510215317,58.6332896898589 21.9845666890459,58.6382493078301 21.9347779264534,58.663448418463 21.8943650901482,58.6914309303908 21.8401040451468,58.7280327803024 21.7990127683807,58.8024397967133 21.7205115184638,58.7950775911053 21.6760432506166,58.802488266457 21.6148680261066,58.8480488999374 21.5935700156607,58.8688836672235 21.5939640265429,58.8859267519012 21.6062946274745,58.8954042203704 21.6187097107752,58.9161844493334 21.658065424624,58.9967498416596 21.6864656094361,59.003217761385 21.8092019608218,59.0080564118485 21.8946637595807,59.0063852256435 21.9605942956779,59.0130992180397 22.0757031128032,59.0340052142756 22.1053510244001,59.0365995639761 22.1214654755141,59.0430958301371 22.126957993053,59.0533764143827 22.1421999900346,59.0417927325163 22.1760867721844,59.0168293845203 22.2071179919954,59.0126037496748 22.2259469977024,59.0118048317269 22.3501207717276,59.0007620171919 22.3612699594903,59.0007021306189 22.3777937487495,59.0034754767876 22.3809426214505,58.9918883004013 22.3875105357664,58.964782559812 22.413483659937,58.9445792584638 22.4302514591467,58.9355697599668 22.4427522576202,58.9374234812086 22.4482378017567,58.9566149780496 22.4607669083376,58.9647240994262 22.4724170222006,58.9661038543778 22.4919330389927,58.9400184361481 22.4856594436245,58.9327796940905 22.4876278075847,58.9262219812774 22.4980493133067,58.919632659396 22.4998507053194,58.8950488757042 22.4911516176065,58.8829370611763 22.4969844794245,58.8832565817897 22.5155068810279,58.889617535733 22.5295289409484,58.9025663090889 22.5469202194522,58.9009016276786 22.5580631274103,58.8847784217128 22.5860071143031,58.8739936650135 22.599902931053,58.8432081602316 22.6266973013434,58.8396583117527 22.6322427399342,58.8395780240146 22.6601301231717,58.841729599172 22.6747802402113))",Wilayat Bidiyah,ولاية بدية
"POLYGON ((58.3760733538487 22.9847765572598,58.3675501567373 22.9866421155164,58.3423127374054 22.9800687616881,58.3316191184677 22.9788873426482,58.3183499759453 22.9638798600236,58.3065854139723 22.9471703544567,58.3049550939641 22.9354491750581,58.3072899418686 22.9244089741349,58.305720413616 22.9111118294891,58.293552454834 22.8913170034678,58.287546142367 22.8914921250943,58.2912732238926 22.8760755458946,58.3017567588461 22.8048638031157,58.2856979410853 22.7716546049589,58.2860712161467 22.760536735809,58.2987238669649 22.7576032147915,58.3217517627791 22.7578500615446,58.3480450907373 22.7556691266888,58.3592720567822 22.7505622158481,58.3668716382378 22.7343655070994,58.366084720615 22.7260919699247,58.3514339771069 22.7101446841845,58.3463654470342 22.7011125129592,58.3466472282369 22.675823061049,58.353881167675 22.6585412028102,58.3548491910013 22.6422296463201,58.3523298415636 22.631780837078,58.3531837790343 22.6202565334187,58.3723627545848 22.6046876788785,58.3794078448284 22.5942165277419,58.361431367417 22.5823089516702,58.358867140042 22.5729182638197,58.3653777189842 22.5688455956304,58.3745297420688 22.5694562908617,58.3847163569436 22.5746489325737,58.3964286094309 22.5753386001599,58.4210431379664 22.5700577617672,58.4338168206208 22.5746634185479,58.4530163897223 22.5661043858932,58.4661677184414 22.5657174338085,58.4894146577752 22.5701623042403,58.5560364801998 22.5783806425982,58.5681486434628 22.5704276958206,58.5927083792676 22.564113376626,58.6002239133616 22.5568303878871,58.6094632432081 22.5588405845308,58.6069879415709 22.5684764401063,58.5899867348593 22.5812796104578,58.5840400854526 22.5902870089286,58.5897173769806 22.5989381902599,58.6171386610115 22.6339316530866,58.61480384898 22.6424329831683,58.6202680824847 22.6515293299689,58.6082226606508 22.6670895181534,58.5865463686422 22.7070301173093,58.5809028182967 22.7097510450978,58.5830114168743 22.7197886134275,58.5741077488173 22.7253388506407,58.5730254416173 22.7369445713559,58.5756001355032 22.7557856389463,58.5754575075161 22.7704064748496,58.5721416671839 22.7761130922031,58.5719609689433 22.7883906639716,58.5797238897254 22.8000681518259,58.5828347399612 22.8104101387205,58.6131164650749 22.8213537507427,58.6255223069169 22.8324202724074,58.6395058226614 22.8332905539742,58.6497226088593 22.8442222660731,58.6585874777142 22.8419756288732,58.6669929057621 22.8465817145854,58.7036104929965 22.8579670015919,58.718843406408 22.8897675770006,58.724694460394 22.9047841648132,58.7233040179018 22.9085869322208,58.709167830712 22.9062355239867,58.6978255670053 22.9078223997699,58.6867408064557 22.9023255898273,58.6799850752812 22.9061968935971,58.6727221899272 22.9025325065768,58.6632897773327 22.9050269801826,58.6554518403269 22.9122184312225,58.6475022188731 22.9128113414371,58.6400575066581 22.9209372253533,58.6271343740227 22.9187695448594,58.6226342227425 22.9216648749318,58.6089372082733 22.9185553492451,58.5982183747665 22.9121092908446,58.5902841619035 22.913638425248,58.5750885516847 22.9114869127554,58.56566065341 22.9144520434017,58.5512153389138 22.9118234670624,58.5412728537718 22.9063005607993,58.5316457417511 22.9205885886174,58.5165129415051 22.9243125002632,58.5088615719203 22.9359161526789,58.4820313871336 22.9376049663842,58.4620456389829 22.9436562825803,58.4544506980851 22.9436877030267,58.4377564117775 22.9506586538215,58.4299074495694 22.9506889591958,58.397511199483 22.9672641692613,58.3760733538487 22.9847765572598))",Wilayat Ibra,ولاية إبراء
"POLYGON ((58.8510008568142 23.363473606533,58.8294695342696 23.3609851028518,58.8254447943019 23.3656283147251,58.804645081404 23.366684601093,58.7997365803019 23.3621403907487,58.7841861356948 23.3739175409875,58.7786089839072 23.3706851116481,58.7671407464236 23.3748831431013,58.7633051984036 23.3866293942441,58.7688223606169 23.3919467081115,58.7642001165184 23.3980603649559,58.7516019737113 23.3892826162763,58.7399596612268 23.3896158196789,58.7280476162445 23.3952766795448,58.7219419329543 23.3918132688624,58.7146580431176 23.3791607395148,58.7156719511141 23.3726704333761,58.7003403999014 23.3673541273732,58.6882046603499 23.3749218574506,58.6919014872797 23.3841083948085,58.6844763513197 23.3868050405027,58.674774732773 23.3797713421399,58.6655325258218 23.3793214619203,58.6623486957117 23.38797710076,58.6720321074424 23.4006291896654,58.6547429977717 23.4133225701908,58.656230209715 23.4258836650048,58.6495079369714 23.4293967135926,58.6345923660847 23.4214363764844,58.6226341876613 23.4118646205401,58.6255631213109 23.4028646495428,58.6172525205831 23.3967785347809,58.6243313918009 23.3902244983827,58.6163729554265 23.384819937205,58.6206066818597 23.375935204278,58.6344148283239 23.3710866482078,58.6414001474914 23.3630197984674,58.638270257022 23.3436420579431,58.664326730758 23.3372300337437,58.6568020714895 23.3267396812778,58.6510082979457 23.3072588722463,58.6486338107098 23.2767904015974,58.6515934640506 23.2599335263041,58.6551410075431 23.2577900360585,58.6570281828067 23.2362084829656,58.6529235647498 23.2294956102664,58.6442717592705 23.2304163790255,58.6376798841718 23.2244911371558,58.641809496159 23.2158519148404,58.6406000435988 23.2047749193978,58.6473923208393 23.1922022590651,58.6411442251497 23.186115638809,58.6499532761094 23.181007638388,58.6756257294649 23.1718062502683,58.6686140790815 23.1547878735037,58.6815602656964 23.1505744036892,58.7275880695939 23.1499790022399,58.7464969231572 23.1480524168837,58.7858179790573 23.1600310502869,58.7919037606343 23.15277881436,58.7910000700562 23.125194597114,58.7958086227328 23.1202734318818,58.8049047693354 23.0636760512512,58.8368641958279 23.045735579718,58.8986916559419 23.0081974511675,58.9118702581573 22.9833644344425,58.9076525564895 22.9658488218295,58.9153821712746 22.959821037656,58.9579629195108 22.9601451985695,58.9664441471785 22.9297611258222,58.9818551919867 22.9150894207549,58.9924621230117 22.8960851919588,58.9821420695898 22.8819715120434,59.0088044388239 22.8720485648484,59.0324104951121 22.8617534562117,59.054795527886 22.8541232872872,59.0766402572923 22.8426246080564,59.1573411833883 22.8411020768918,59.2248222981229 22.8852911997083,59.2252129284738 22.8963622175979,59.2177962600384 22.9162290779711,59.2126895818738 22.9235990438593,59.2063601324139 22.9436771580454,59.1959965178618 22.9585377396712,59.1830123053773 22.9702307069485,59.1603371501466 22.9785439101454,59.1420938995865 22.9917329482384,59.1209692433508 23.0005587360102,59.1050295068168 23.012620644014,59.0938352929917 23.0247645420637,59.073958917179 23.0413006519713,59.0655508924038 23.0540277155746,59.0584884328657 23.0816604994242,59.045866749714 23.0929030859626,59.02819776382 23.1035419192248,59.0138179436297 23.1194994459895,58.9980842908468 23.14637836683,58.9898114797062 23.1714684238987,58.9939554519412 23.1890446630348,58.9887882476098 23.2081177881904,58.9587709058529 23.2330712902986,58.9429151315657 23.2396401508077,58.9248558050791 23.2592204654102,58.9261804066724 23.2680649754154,58.9204202741065 23.2777841787408,58.917120828733 23.3013048126903,58.9083762814922 23.323727683821,58.8954660299491 23.3262739511164,58.8830856473342 23.334933603293,58.8761100713649 23.3451144687891,58.8667417296446 23.348772915469,58.8510008568142 23.363473606533))",Wilayat Qurayyat,ولاية قريات
"MULTIPOLYGON (((59.8232483508265 22.360452949277,59.8234470818067 22.3679393365161,59.8168419538806 22.3780315086213,59.8182465543987 22.3909938435541,59.8297524891871 22.4174417347658,59.8377867969285 22.4229822189901,59.8372982173425 22.4315452838047,59.8247269511828 22.47446046433,59.8156909792993 22.4924872461283,59.8078225941473 22.4980592442569,59.7952677959426 22.5381328239667,59.7842189139521 22.5383584946086,59.7622656368574 22.5321245481336,59.7662354149978 22.5279953002555,59.7840058751382 22.5263231901576,59.7851229592496 22.5179526641214,59.7603044998707 22.519751207167,59.7611292258876 22.5244203174254,59.7529510013624 22.5331322963702,59.7355727320537 22.5357173192038,59.7340864537211 22.5295449112944,59.7287430030404 22.5258111142711,59.7391562162552 22.5147758098409,59.7507944249021 22.4976879062862,59.7630880015662 22.4959685563905,59.7651612154607 22.4890139773384,59.7551471458369 22.4836608880362,59.739214768719 22.4820632602987,59.7244793955602 22.4954061080979,59.7145085195271 22.4999979204953,59.7138860556448 22.5070105760727,59.7258564177999 22.5171025529146,59.7291961262899 22.5231316745894,59.7267879432907 22.5249855882213,59.7307643973219 22.5276663730399,59.7319850778024 22.5343667289388,59.7282074085574 22.5372808854244,59.6982669711709 22.5422733183336,59.6714984621396 22.5525394487361,59.6487469485749 22.5590269186414,59.6365645976992 22.5586327453687,59.5951525678736 22.5630479311739,59.5925442808725 22.5655417900146,59.5596393937965 22.5664838677786,59.5420073959375 22.5695432905708,59.5363221004489 22.5536656841285,59.5141817542182 22.5501651603518,59.5102532220927 22.5574292145482,59.5124215419152 22.5677787636545,59.5218730374672 22.5616151301095,59.5361469455567 22.5599349368055,59.5379166692992 22.5674724294579,59.5288841012721 22.5756356902126,59.5033658661761 22.5917239724557,59.4855290544617 22.6015126525782,59.4616800187243 22.6181230248881,59.4227215628558 22.6556339326364,59.401330980412 22.666971504114,59.3832404403635 22.6811079038244,59.3762060225472 22.7060504814552,59.3582839977152 22.7099426289528,59.3488778052154 22.7228529100624,59.3410954308031 22.7438642311984,59.3346600815031 22.7518582046407,59.3188108208556 22.7568519341188,59.3053639190132 22.755564469261,59.2926919280031 22.763039930229,59.2835743803483 22.7764352721486,59.281440111898 22.7862680671494,59.2653998266187 22.8144347171867,59.2638710630982 22.8248316808091,59.2571864419278 22.8294661494649,59.2407943998847 22.8471008124656,59.2341981297122 22.8697406819167,59.2248222981229 22.8852911997083,59.1573411833883 22.8411020768918,59.0766402572923 22.8426246080564,59.054795527886 22.8541232872872,59.0324104951121 22.8617534562117,59.0088044388239 22.8720485648484,59.0136686918132 22.8605868838761,59.0228794873163 22.8503455237104,59.0430700319762 22.8341503607002,59.0474775363124 22.8254050282738,59.0666613859709 22.8186085958939,59.067280096738 22.8069276561337,59.0749994832871 22.7962075389859,59.0874498589347 22.7852846720839,59.0909659444005 22.7752958246149,59.0899181080606 22.7528074085357,59.0913527776265 22.7472541781927,59.1007777674698 22.7329208301466,59.1185539223589 22.7171159238787,59.1242942632743 22.7052476423795,59.151233219355 22.6786170055577,59.1406205141571 22.6715561222059,59.1376989123511 22.6611030236993,59.1527862499431 22.6390161007814,59.170037231398 22.6253727384013,59.1799654047164 22.610423341405,59.1930619181616 22.6045835459762,59.205755722366 22.5869336299465,59.2055832542139 22.5682794689524,59.1969960072709 22.5620179758383,59.1977265535305 22.5519494280398,59.2076638763575 22.5439759285805,59.2134668727311 22.5451534667415,59.2149444462081 22.5311875658368,59.2199517431622 22.5192158544764,59.2331441681103 22.5035754938877,59.2484920064373 22.4953034792113,59.2539131847511 22.4970177183618,59.2590362810292 22.4811541803344,59.279635769476 22.4599665915565,59.2915917184511 22.4568108319012,59.3038829206835 22.4403657172698,59.3246002191719 22.421586697767,59.3621676585898 22.4052806311723,59.3652619442479 22.3934340457156,59.363677211843 22.385906560427,59.3735038181256 22.3676066071158,59.3817720073295 22.3571270516784,59.3978379964327 22.3450805164122,59.4051327308771 22.3443628964766,59.4192415029776 22.3481635810561,59.42192239865 22.3588808371624,59.4292494145712 22.3652736923223,59.4463907405527 22.3711975231957,59.454274869822 22.3602735525023,59.4685299698081 22.3680940471434,59.4759486594778 22.3665677727163,59.4875470243662 22.3710483367528,59.5041278906553 22.3644909618743,59.5135826083804 22.3681812260475,59.5173877139838 22.3741910783058,59.522260247519 22.3942857194129,59.5358171966832 22.416889168649,59.5450109484815 22.4251524009108,59.5622919408316 22.4260255689457,59.6181154114187 22.4216904674893,59.6540143480354 22.40734689121,59.6799520152513 22.399235125303,59.6942466208153 22.3646565192907,59.704631130374 22.3677845673031,59.7135054691501 22.3553767751266,59.7916656907279 22.3605174280422,59.8232483508265 22.360452949277)),((59.7133277186826 22.2779290011056,59.6955544648458 22.2705691655549,59.690184334102 22.2645247250681,59.6756702559208 22.2622570500416,59.6816733800669 22.2473544630944,59.6867521258682 22.243186204368,59.6932525817998 22.2502908738251,59.7037200790295 22.2407988114637,59.7055466821681 22.2346105308068,59.7159290028346 22.2383312845649,59.733743193385 22.2390286729475,59.7358872356286 22.2442447961554,59.7288471992103 22.251564918983,59.7224363943284 22.2768438444484,59.7133277186826 22.2779290011056)))",Wilayat Sur,ولاية صور
"MULTIPOLYGON (((57.058891250751 24.0224231987734,57.0462707406998 24.0121700110424,57.020981315412 24.0337904790356,56.9969828300034 24.0444363236558,56.9839253396404 24.0294505330206,56.9667911376202 24.0212096858126,56.8969042991333 23.9717925220927,56.8963226418863 23.9667527877276,56.8826860868881 23.9527476365771,56.8716274186591 23.9191181815662,56.8614418462245 23.8940758614896,56.9381574569653 23.893084118321,56.9485052787326 23.8728271202045,56.9153337080125 23.8016187266885,56.9077360266087 23.7666250903258,56.8998612324199 23.7232471551562,56.8993728424919 23.7137135523303,56.8901362341169 23.6839336254225,56.8927118544688 23.6163858174042,56.8848922287047 23.5964730407166,56.9184561766945 23.5904156845971,56.9172358517373 23.5575858518087,56.9255450165945 23.5443881516878,56.9485447722418 23.5317235001861,56.959710611883 23.5333182228394,56.9866105451378 23.5412368579328,57.0041785903287 23.5635385770995,57.0360308316768 23.547668422976,57.0909877707499 23.5647534226562,57.0416869804616 23.6308093871864,57.0454157095675 23.655791147101,57.0753594287983 23.6607331869273,57.1030783076364 23.6987133594241,57.1316368904858 23.7603178491982,57.139077669174 23.7813307715453,57.1609345582231 23.8092907268387,57.1631038455383 23.8209689799977,57.1606781928452 23.8274683318758,57.129809038168 23.8544390712902,57.1188784905335 23.8698430908918,57.1201831909695 23.8881978461004,57.1296629295869 23.8976201136269,57.1474968880666 23.9355898620164,57.1578851129231 23.9470759055079,57.1397119036886 23.9575439416742,57.1207888211262 23.970977132187,57.0985661762121 23.9893965209832,57.0798281228615 24.0082713664027,57.058891250751 24.0224231987734)),((56.5498596450383 23.7831032543773,56.5606638530844 23.7785523401547,56.5701032325482 23.778289873231,56.6321682161665 23.8031143046281,56.6539332483305 23.7875218495692,56.6401329881716 23.769023072177,56.6477307172913 23.7528183475121,56.6926186893222 23.7353882562129,56.7114142195637 23.7896935502149,56.7226791319721 23.786683712279,56.7291382683574 23.7785679591413,56.7358414397874 23.7768046582167,56.7772425792622 23.7905373796658,56.8260396159744 23.8450922992754,56.8045857476312 23.8747226205568,56.8228981109326 23.922873171815,56.7803443402806 23.9674135421636,56.7747578380811 23.9680022600898,56.7355672040349 23.9598981000461,56.723218540988 23.9764822427098,56.6910543491704 23.9839155317281,56.6651997178926 23.9622883901113,56.6559944887482 23.9359631618412,56.6467273946181 23.92198140935,56.5979965056291 23.9061620473095,56.590887479378 23.8849406042133,56.5785864136235 23.8814640597083,56.5718119449887 23.8533327625855,56.518024239392 23.8318598840931,56.5411386378796 23.8173927328728,56.5498596450383 23.7831032543773)))",Wilayat Al Khaburah,ولاية الخابورة
"POLYGON ((57.4665875616156 20.989135143368,57.3391767426874 21.0115322059444,57.1221718176992 21.0599769344571,56.7075739395412 21.2359829222017,56.6861257076206 21.2212003416346,56.6518802274495 21.2298853091513,56.6315664404592 21.2655798309765,56.6288489946401 21.2730143513206,56.5262051183743 21.3277858407854,56.577367899338 21.4908794452847,55.4439124493263 21.3373088530363,54.9999999983451 20.0000000436826,55.0102061953275 19.9845643688199,55.0573749325999 19.9984070021751,55.0874155273192 19.961681388719,55.0553759604434 19.9162032802052,55.6891378079147 18.9490818683714,55.8402280132996 18.7163673047502,55.9186973266928 18.7566464331016,55.9655442654266 18.7877119814003,56.004876752186 18.7991482680057,56.0180136869433 18.7992392998394,56.0509643973851 18.7910061213276,56.0789019530524 18.7857850809901,56.1273847805011 18.7833368111428,56.1269270736877 18.8719792241844,56.0978320989593 18.9028226016464,56.0777085363308 18.9448936318646,56.079446577496 18.9578113732898,56.0784617047 18.9724367643168,56.0852670095965 19.0044544104995,56.1015368152674 19.0551682353469,56.0916147462422 19.0883767890257,56.1095068726772 19.1172814538915,56.1469182002006 19.1178751056816,56.1572334900845 19.1053461727701,56.159302034385 19.0947780549616,56.1940951797382 19.0379639728825,56.2475812029582 18.9853836513755,56.3000658008617 18.9785705896532,56.3015591597526 18.9793905976889,56.4002399026315 19.0816387684353,56.4122801833183 19.0945469181164,56.4282124695064 19.1010317462257,56.4393388448401 19.0992274675466,56.455891366393 19.090465138602,56.4705965934749 19.0950268283152,56.4865396656246 19.0938157204497,56.5854881638252 19.1607582717855,56.6025411008747 19.1751300734416,56.648537834905 19.2059916058296,56.7494202008881 19.245426996549,56.8031912498422 19.2567397602619,56.8635382327898 19.2792413821969,56.9864847450524 19.3185977099406,57.0446862435819 19.335409009436,57.0787347402994 19.3438293261446,57.0897178017582 19.3494386952711,57.1113161180224 19.3727014418215,57.2497924664554 19.5538467721999,57.3060555323464 19.7603461621647,57.3285178410388 19.7841044811833,57.339894335995 19.8585859349464,57.3926162757057 19.8974519376903,57.4049842306293 19.9207390298585,57.3961588160557 19.9429048861478,57.3710493243599 19.9360787750025,57.3595976467853 19.9297399709134,57.34143733598 19.9316844946072,57.3267392886675 19.9816565419022,57.2864687898224 20.0415320276561,57.2807517732975 20.055709923789,57.2832083474687 20.1477186457019,57.2935710745365 20.1725990329458,57.2936258157997 20.2018261841141,57.3349347404539 20.2158246142155,57.3865456472626 20.2189660484392,57.399231750539 20.2470820360565,57.3889657664219 20.2698370422906,57.3718027496603 20.2882763320065,57.348961776509 20.3348695709239,57.3581700655025 20.3467580736534,57.3616509424294 20.3629878688884,57.3536458316756 20.3759938170831,57.3387229683337 20.3760234209214,57.3330019943814 20.3846941437157,57.3491297490045 20.4095591949979,57.3744416002119 20.4311557472657,57.3894324162231 20.4560192258095,57.3940982408966 20.4841523378482,57.4067711437722 20.4981948914322,57.4033615326527 20.5122745775466,57.44243704029 20.516509110218,57.4562756720392 20.5337922054144,57.4551874724619 20.5543612608534,57.4518225787715 20.5825132130925,57.4565040859986 20.6106439685752,57.4450548030627 20.6269101683123,57.4232271138168 20.6334595665404,57.3656944622002 20.6162720730519,57.338163768365 20.6444713676961,57.3658887163988 20.6974536381442,57.4108353044952 20.7287423493979,57.4328279740097 20.7752319654679,57.5156841077731 20.772838385412,57.5284263926757 20.7966122859438,57.5227234289762 20.8117832204638,57.5077765667836 20.817240084704,57.4502551077049 20.830389544455,57.4688672051316 20.8920358676656,57.4758836646696 20.9255703584454,57.4682687699987 20.9611358979306,57.4665875616156 20.989135143368))",Wilayat Hayma,ولاية هيماء
"POLYGON ((56.2869242156172 25.3294767491741,56.2760322338546 25.3372974508149,56.2657149333357 25.3343817330345,56.2480610726453 25.3249089630658,56.2440247727287 25.3170629226477,56.2586042807977 25.2964023817598,56.2553598190181 25.2823915848732,56.246881562806 25.2818916226411,56.2379546238767 25.2727636211252,56.2233846975022 25.2622119667089,56.2244248056964 25.2487826786515,56.2342787377955 25.2478745401962,56.2475545238778 25.2405376587724,56.2583936567512 25.2378640513304,56.2606561761162 25.2430647539755,56.2721293449904 25.2425866874157,56.2821636600627 25.2366975259921,56.3049406870914 25.257862630156,56.3213182056666 25.2611845135176,56.3377626965175 25.2729238253524,56.3448813403876 25.2743932320266,56.350575617431 25.3042897742878,56.348957593944 25.3064957970054,56.3226502159682 25.3098733780466,56.3197399201821 25.3024527742823,56.3092732274746 25.3152937835193,56.3096853421071 25.3218280420073,56.3032866418281 25.3298467017046,56.2910563916716 25.3251807695819,56.2869242156172 25.3294767491741),(56.2691875216968 25.2821310270003,56.2777857813916 25.2903814413701,56.2890772126085 25.2754045394841,56.2846375321984 25.2627741479435,56.2700025481908 25.2640871232647,56.2691875216968 25.2821310270003))",Wilayat Madha,ولاية مدحاء
"POLYGON ((56.8414913653767 24.2393476107999,56.8296907735265 24.2533572339234,56.7689924954685 24.3395385039893,56.7356111089042 24.3831851749223,56.7187970857628 24.4093207716431,56.6930242807557 24.4248980433075,56.6514669154304 24.4613571426938,56.6309847876482 24.4816747447056,56.6315581623242 24.4890734447653,56.6032418590528 24.5227586929542,56.5837918629657 24.5114456638156,56.6211558116319 24.454402267734,56.6102078880428 24.4486008667109,56.5705506861093 24.4529307949604,56.5662591564109 24.451680106998,56.5594766838877 24.4388237198414,56.5427574436415 24.4315782992542,56.5344352864255 24.4179434524981,56.5339710064081 24.4048018244358,56.529574454122 24.3967020543107,56.4944876706013 24.3867425859019,56.4731402791766 24.3855327262649,56.4390051969048 24.3626835335924,56.4362030431712 24.3343753773861,56.4108570786259 24.3352569906318,56.40311480564 24.322518259343,56.3899489261408 24.318397323314,56.3866174562856 24.3117261954428,56.3667127733963 24.3104115843376,56.3607000680146 24.3290032358267,56.3526380889385 24.3372659420121,56.3260715090555 24.3381752190403,56.280900203305 24.3108876127464,56.2807093972695 24.2794860850053,56.2915857356622 24.2416946448008,56.2799106579318 24.2340067593173,56.2776358577937 24.2218477478202,56.291851716719 24.2148189599381,56.2961834668668 24.2026491162786,56.2747455488995 24.187616859336,56.3002526652494 24.1781974172092,56.3010169449498 24.1669125538614,56.3122820884177 24.162770903461,56.3368422332675 24.1465382287356,56.342985018495 24.1360287468725,56.3457616124799 24.1195916991177,56.3518904267381 24.1114470592511,56.3492649359882 24.0982121185531,56.3539300215701 24.0918487211834,56.3580958476392 24.0642761173073,56.3680290169707 24.0192702024349,56.3923618332818 24.0191536627525,56.3995604981715 24.0056354834704,56.4038986998768 24.0033946055974,56.4021805932562 23.9920978763402,56.3801462113188 23.9854300001745,56.366095289422 23.9764176849778,56.3773207647941 23.9744963081262,56.3903805601555 23.9590132852871,56.3954714206649 23.9590334154566,56.3970739512362 23.9471403379448,56.4014576689634 23.9398592916329,56.3832749616439 23.9301834479269,56.4062985821457 23.9139597283266,56.4393659729854 23.9160925606266,56.4606808425383 23.9090062207439,56.4663178334335 23.9012920328476,56.4741337093871 23.9016581108768,56.4854548428578 23.8921986298928,56.4842043452951 23.8727917874405,56.4926251315816 23.8688848934993,56.4959760999532 23.8603478151807,56.4937435796985 23.8467042771889,56.518024239392 23.8318598840931,56.5718119449887 23.8533327625855,56.5785864136235 23.8814640597083,56.590887479378 23.8849406042133,56.5979965056291 23.9061620473095,56.6467273946181 23.92198140935,56.6559944887482 23.9359631618412,56.6093817907965 23.9872646680539,56.5556043910468 24.0077093546925,56.5596722686423 24.0105396001834,56.5717893424014 24.0392790543121,56.5864121953945 24.0385411519884,56.592306437568 24.0540718132166,56.6036011852927 24.0940778989977,56.6693598797609 24.1790418303609,56.7864522319653 24.210763587348,56.8093952838272 24.2238310256967,56.816861202911 24.2313942084522,56.8302897859773 24.2283450130693,56.8414913653767 24.2393476107999))",Wilayat Sohar,ولاية صحار
"MULTIPOLYGON (((58.8908380092862 20.6963263319196,58.8722346896647 20.6900088196493,58.876330087964 20.6767227953895,58.8714567470456 20.6624748786474,58.8712033569043 20.6527221804635,58.8632770529737 20.6365687466923,58.865337299439 20.6176573319299,58.8406566000207 20.6019033736406,58.8256311899699 20.5839336869431,58.8178943064494 20.5718854561108,58.811492404943 20.5557361832841,58.8063575060046 20.5522614043853,58.7857062323611 20.5202421775046,58.7853556147767 20.5019418196336,58.7810996313066 20.4808982674565,58.7845000735301 20.4714159214761,58.7778329828783 20.4618882222753,58.7740495767117 20.4414390485751,58.7677089204976 20.4339956464366,58.7573763746144 20.4305431012094,58.7514182226006 20.4224592503357,58.7339695655683 20.4239524112522,58.724656116821 20.4211499445548,58.7171586193347 20.4298962749944,58.7048020547831 20.4287834540465,58.6991697116666 20.4168765169885,58.689253076711 20.4134319180852,58.6843581795661 20.4072926560917,58.6827094329609 20.3921314535099,58.658839079553 20.3776795069041,58.6522903856675 20.3698018872562,58.6381736183123 20.3467852972364,58.6330760997096 20.3447044397363,58.6314998979884 20.3233010550799,58.6340234119476 20.311306151108,58.6325348897135 20.2965440140945,58.6234282261895 20.2695423924605,58.6288426765376 20.246631721961,58.625270675201 20.2386713806827,58.6266440074504 20.2248937461804,58.6348537755787 20.2162196266547,58.6343933207055 20.19578080651,58.6294276431483 20.1863433211221,58.6342633118051 20.1803821306067,58.6341038583203 20.1717899777167,58.6447645869749 20.1683951692768,58.6585714797415 20.1691270099449,58.6668098459976 20.1858316431108,58.6717854698247 20.1898952033705,58.6909823705121 20.1970044397693,58.7136758575511 20.209593360816,58.7235077150537 20.2169333545738,58.7332116326538 20.2393444353748,58.7388907010375 20.2483044222686,58.7682270050971 20.2692216010719,58.7820502577195 20.2776528938456,58.7778666100979 20.2835536407362,58.7776676754195 20.3000203743226,58.7935091806208 20.3212674735575,58.8010560938226 20.3555497413238,58.7981617221447 20.3599987204926,58.816466035385 20.3849133296053,58.8209731804503 20.3964771572804,58.8187717827662 20.4071970026481,58.8234889270241 20.4186252834797,58.8466909669681 20.4445739886381,58.8879957390455 20.468045845878,58.9041893813491 20.4741218030413,58.9049466232898 20.4792122137902,58.9161870800116 20.4852210882148,58.9281974550463 20.4876497914448,58.946685356274 20.4957667869334,58.9510460387877 20.5049092511333,58.9610475109966 20.5153841770995,58.9584364467616 20.5206067885706,58.9464822837042 20.5242725135095,58.9371613599058 20.5418722277176,58.9382892203091 20.551658813797,58.9351336540508 20.5603245722787,58.9377540537026 20.5735513782248,58.9124336816431 20.5873824138964,58.9085887044469 20.592946351255,58.9008024375486 20.6174390679468,58.90089417948 20.6254381649995,58.9076160759528 20.6560684134377,58.9127175417724 20.6666935409648,58.9148376346308 20.6855475425087,58.9116628126308 20.6923492990469,58.8908380092862 20.6963263319196)),((58.7512476266143 20.4722977419701,58.7464914832433 20.4727395157543,58.7418701023818 20.4617741526815,58.7403978283381 20.4490105758807,58.7531754307456 20.4547249516529,58.7572277156715 20.4619231728228,58.7512476266143 20.4722977419701)))",Wilayat Masirah,ولاية مصيرة
"POLYGON ((57.6951789063901 23.1562320103669,57.6745225981536 23.1516538592947,57.6254189111624 23.155427904989,57.6148477758737 23.1610017117779,57.6053570126213 23.1545259142653,57.5932300375817 23.1679473606814,57.5411958732754 23.1793392438928,57.5043366156789 23.1817025339094,57.4976552966017 23.164894661691,57.4632023306488 23.1509576653776,57.4429423167376 23.1553541340959,57.4378052262602 23.1516051941218,57.4297181418011 23.1084945415168,57.4069350089254 23.0784414025226,57.3896902552256 23.0737021289662,57.3649928516505 23.0735839693801,57.3418177695608 23.0492355567763,57.3372691882338 23.0484531624246,57.3438195317748 23.0358462140596,57.3541188158461 23.0327868855031,57.3549300313934 23.0247897907957,57.3669994475878 23.0110875801297,57.4058890848277 23.0078882326807,57.4218334497852 22.9485395908336,57.3844328308752 22.9189007658775,57.3784251361324 22.8697678743613,57.390910948859 22.8511961329099,57.3797556213022 22.7723591745184,57.4789929840942 22.6862691275745,57.5290406914977 22.7482457803368,57.5554875179866 22.7780673765756,57.5648640386637 22.8283951376657,57.5999156353851 22.8302290877283,57.6291797833739 22.8571056698022,57.6572502949887 22.8731247677458,57.6963889938017 22.8772161150716,57.732812946825 22.8845917339745,57.7251716134998 22.9241789278708,57.7263447325872 22.9388771366702,57.6969033549002 22.9608448764559,57.7131896224724 22.98712305299,57.7368914189014 23.0069873825142,57.8066596186993 23.0904063239876,57.7873093976885 23.1426732898508,57.7574451686242 23.1193450072182,57.7351207964276 23.1189604059127,57.7194516355502 23.1320575903342,57.7209750331172 23.1621620425334,57.6951789063901 23.1562320103669))",Wilayat Nizwa,ولاية نزوى
"MULTIPOLYGON (((56.366095289422 23.9764176849778,56.3801462113188 23.9854300001745,56.4021805932562 23.9920978763402,56.4038986998768 24.0033946055974,56.3995604981715 24.0056354834704,56.3923618332818 24.0191536627525,56.3680290169707 24.0192702024349,56.3580958476392 24.0642761173073,56.3539300215701 24.0918487211834,56.3492649359882 24.0982121185531,56.3518904267381 24.1114470592511,56.3457616124799 24.1195916991177,56.342985018495 24.1360287468725,56.3368422332675 24.1465382287356,56.3122820884177 24.162770903461,56.3010169449498 24.1669125538614,56.3002526652494 24.1781974172092,56.2747455488995 24.187616859336,56.2961834668668 24.2026491162786,56.291851716719 24.2148189599381,56.2776358577937 24.2218477478202,56.2799106579318 24.2340067593173,56.2470283805866 24.2318563247062,56.1863863386403 24.2067461890657,56.1522743185627 24.1985564538884,56.1423241792752 24.1868487347807,56.1453659820588 24.1670199635455,56.1429153523436 24.1627413515873,56.1211765474498 24.156840154174,56.1398343366645 24.1083155072379,56.1012159671884 24.0937699670105,56.0622363517928 24.0728920588587,56.0607040207439 24.0641682708158,56.0479139687994 24.0651352585753,56.038114346277 24.0722049608876,56.0178146694083 24.0674136342376,55.9917632941775 24.0628363648929,55.9598733944511 24.060527136087,55.9416463540679 24.0544263185418,55.8990427253249 24.0451132002509,55.8548689606509 24.0219879740725,55.8429336736135 24.0206472337413,55.8337444061063 24.0137484946722,55.8197564968778 24.0208511950855,55.8018622956106 24.0250079598195,55.7801649339402 24.0552890708394,55.7583501544369 24.051312220544,55.74323273257 24.0570128722721,55.7267899970408 24.0555296055929,55.7810220304417 23.963387457889,55.7954421984804 23.9616810570966,55.8206201634311 23.9551819780151,55.8508339233015 23.9551132189633,55.8697781698017 23.9256990488003,55.9017981907999 23.9516539138366,55.9145414672204 23.9153413168619,55.9191724432287 23.8209455096804,55.9556576564907 23.8254409836056,55.9583505844873 23.7867846646571,56.001553811727 23.7843136991836,56.0050295125467 23.8070601784067,56.0008001893264 23.8456139100185,55.9612248017993 23.8986878881513,56.0443963640888 23.9422538863052,56.0689328201332 23.9465518998928,56.0688203279901 23.9622188486238,56.0626717479292 23.9742479129458,56.0491477429145 24.0150770941752,56.1763086486729 24.0135549421218,56.232149805596 23.9817689174369,56.2952571303968 23.9737116853177,56.3450448348159 23.9724893199336,56.366095289422 23.9764176849778)),((55.9472184857905 24.2224983515952,55.9424360869097 24.2308079407951,55.8679265976322 24.3203618128097,55.8299604002969 24.3245630827451,55.8079838309078 24.3104191127504,55.7915958494256 24.2793476682228,55.7679249135996 24.2621803248742,55.7594684971729 24.2610669189347,55.7539346435265 24.2462815382724,55.753003405465 24.2348846366074,55.7656743006224 24.2322688088189,55.7768273570349 24.2348572615922,55.8082040522347 24.2121514618029,55.8138484805151 24.2113662319586,55.8334077505057 24.2013492596425,55.8534235746214 24.211311040896,55.8707650192865 24.2154810069519,55.9472184857905 24.2224983515952)))",Wilayat Al Buraymi,ولاية البريمي
"POLYGON ((53.2273317908702 17.4086275548016,53.1883792625443 17.3827702062217,53.1757628030639 17.3759322643165,53.1708558277822 17.3691737253947,53.1570063390376 17.3676958217968,53.1493623994071 17.3711835447282,53.1409096324381 17.3831370235225,53.1362528475868 17.3945577211089,53.1359852959352 17.4072750634862,53.1438801057085 17.4219681978746,53.1587031772243 17.4374010060192,53.187019694369 17.4482122210308,53.1866057968622 17.468078433119,53.13873965963 17.510436914113,53.1052157204988 17.549854873121,53.0877830999771 17.5920796728692,53.0921941195988 17.5960836239516,53.0918866602642 17.6172407249011,53.0989887983042 17.6347072840721,53.0934330603625 17.6661588143249,53.0832410540031 17.6882894267513,53.0728240445654 17.6895849028656,53.043965042266 17.6978987426785,53.0419947628093 17.7147352383439,53.0200898319925 17.7196256607608,53.0131563609995 17.7322392695085,53.0351258915459 17.7418967033466,53.0495145332738 17.7422752050237,53.0586426459524 17.7726459486622,53.0601359284356 17.8179966629723,53.0373745787168 17.8380991038042,53.035491824974 17.903043171822,53.0586941083733 17.9449813861158,53.056238075992 17.9674185133832,53.0608885107734 17.983337389818,53.0804220551131 17.9953940255254,53.0816047759337 18.0206123531318,53.0815653478731 18.0518442107512,53.0888721914108 18.0757293811523,53.1061469315797 18.1116850638238,53.1352993254534 18.1128974098772,53.1485757690599 18.1231586341157,53.1716091983395 18.1554783499491,53.1786469516003 18.158622745698,53.0059225643277 18.4250246465511,52.6178205315456 19.2107400398903,52.328376689063 19.1123134912328,51.9999999441718 18.9999999600252,52.1957426702874 18.5911880905167,52.782175979986 17.3497337564071,52.7505555123212 17.3058333411362,52.742638813579 17.3019249811302,52.7458333657592 17.2944444708508,52.8122830413653 17.2855303964539,52.9312140511644 17.0315820202588,52.9556181508384 17.0440206774112,52.9713407133697 17.0563730253695,52.9785783347004 17.0427202950107,52.9848986768095 17.0494736672034,52.9932001725295 17.0380795711503,53.0078485957727 17.0459032502182,53.0183727750384 17.0571567004668,53.0640423804939 17.084244191464,53.0802192819321 17.0686276714408,53.0792020039142 17.061258553768,53.0882727455551 17.0492496597762,53.0915497305682 17.0400980040064,53.1046556792866 17.0289934312105,53.1058659581611 17.0152658037964,53.113130439955 16.9965654271656,53.1239136777458 16.990189451488,53.1479778105568 16.9698258965728,53.1572907952285 16.9486013154213,53.1665697012403 16.943009344607,53.1600182558074 16.9360029555175,53.158615811766 16.9251753342951,53.1882110884165 16.9357962434572,53.2469410611709 16.9612614614385,53.2863539249682 16.9872160998117,53.2967628270739 16.9926640418376,53.3644639309539 17.0180045659715,53.3683369426613 17.0325277989031,53.380195213511 17.0468579678559,53.3900912448685 17.0553920767484,53.395772246996 17.0691296022924,53.3987223837785 17.0852185775127,53.3863486983556 17.0921163294725,53.2686730685468 17.0606508409238,53.2547937632091 17.0741294093557,53.2450736402505 17.0760981770581,53.2353291116219 17.0700084981895,53.2272443918922 17.0739763719769,53.2309507161942 17.0840723998219,53.2263363555172 17.0913276566611,53.2176470902304 17.0883006386535,53.2103622673934 17.0802861662393,53.1978939738508 17.080052477889,53.1917632611792 17.0702687142757,53.1826454679482 17.0792285036201,53.1839116355479 17.1084368817402,53.1795175759783 17.1139043140689,53.1660985384993 17.1145455017203,53.1600213763604 17.1203385364834,53.1510432305561 17.1223162281547,53.1300633487249 17.1194090335353,53.1165477449184 17.124699846487,53.1010574209602 17.1442739914299,53.0946138491382 17.1674232965725,53.0853267482288 17.1751204151322,53.0763327439646 17.1734543289349,53.0575714515191 17.175188167068,53.043100939669 17.1806043563941,53.0205831337837 17.1828606718376,52.999074496676 17.1962335099226,52.984843095415 17.2193479123482,52.9745924827323 17.2525853197983,53.2565313718648 17.3658641644997,53.2273317908702 17.4086275548016))",Wilayat Al Mazyunah,ولاية المزيونة
"POLYGON ((53.158615811766 16.9251753342951,53.1600182558074 16.9360029555175,53.1665697012403 16.943009344607,53.1572907952285 16.9486013154213,53.1479778105568 16.9698258965728,53.1239136777458 16.990189451488,53.113130439955 16.9965654271656,53.1058659581611 17.0152658037964,53.1046556792866 17.0289934312105,53.0915497305682 17.0400980040064,53.0882727455551 17.0492496597762,53.0792020039142 17.061258553768,53.0802192819321 17.0686276714408,53.0640423804939 17.084244191464,53.0183727750384 17.0571567004668,53.0078485957727 17.0459032502182,52.9932001725295 17.0380795711503,52.9848986768095 17.0494736672034,52.9785783347004 17.0427202950107,52.9713407133697 17.0563730253695,52.9556181508384 17.0440206774112,52.9312140511644 17.0315820202588,53.1064780701571 16.655581029791,53.1173926542497 16.6531817630919,53.1327477875054 16.6630005012444,53.1508719319159 16.6678733381266,53.1628181722363 16.6770953777088,53.1759554509917 16.6797380461679,53.1895133766388 16.6899131855252,53.2332264417806 16.7011355433765,53.2520686447824 16.704632198651,53.2633662131156 16.7102008872178,53.2929615354538 16.7185768568544,53.3065307600546 16.7189465021155,53.3255695228885 16.7232682230695,53.3317516302658 16.7285408920301,53.3437836172894 16.7317155527608,53.3697443313465 16.7352525259336,53.3474101380974 16.7423641283029,53.3390071658156 16.7388941275927,53.3320287901747 16.7427689590379,53.3162522784802 16.7411464199788,53.3080543225579 16.7468766614933,53.2907972143687 16.7493393703598,53.2651629915255 16.7500730986324,53.2592756080982 16.74821459022,53.2474508804875 16.7567061432602,53.2381844323294 16.754214707265,53.2036950623923 16.7556370018996,53.1935880039937 16.76129287995,53.1846195089798 16.7590843256964,53.1670519524728 16.7602795663432,53.1526103911524 16.7651159444561,53.1358036418982 16.7794762658421,53.1371541810432 16.7901437242966,53.1327604006038 16.823481902673,53.1295177539663 16.8610189642566,53.1380225074517 16.8974555042951,53.1471880142713 16.9142006024052,53.1437558398788 16.9208316662268,53.158615811766 16.9251753342951))",Wilayat Dalkut,ولاية ضلكوت
"POLYGON ((53.754728287116 16.8702802043016,53.7262980225754 16.8686309072435,53.7165402858676 16.8661705217009,53.7109406835001 16.8568898738238,53.6952491214712 16.858683228321,53.683248121309 16.8562472728582,53.6734383125188 16.8492661950838,53.6708331838852 16.8609013392954,53.6564796959297 16.8704131799345,53.6761963476368 16.8924359745873,53.6633331670425 16.9016043146425,53.6582876045839 16.8968268642282,53.6438515273 16.8995760556567,53.6346753997748 16.9041912945753,53.6333551415038 16.919353394597,53.6370160895435 16.9338178941847,53.6295993859583 16.9397038589341,53.6387264587191 16.9521723283728,53.6355512537697 16.9796103774612,53.6284339281638 16.9900028985101,53.6219755591281 16.9926511353509,53.6191106313397 17.0039700792525,53.6061117861869 17.0240966307484,53.596179727064 17.028716634879,53.5890691419138 17.0400820222974,53.5753665704764 17.0424835473781,53.5560626828722 17.0575223938428,53.5539966727127 17.0659061858331,53.5405508885394 17.0720358365901,53.5351339788958 17.0845453992073,53.5352838988151 17.0962152912083,53.5210391787585 17.0925045075454,53.5117323727005 17.0957605466219,53.4812088221007 17.0966388418502,53.4674927155617 17.0899194586136,53.4561024415356 17.0983609212707,53.4475535129536 17.1001702107989,53.4223692432505 17.0977673942284,53.4086168768171 17.09852848514,53.4043229838116 17.0882046656859,53.3987223837785 17.0852185775127,53.395772246996 17.0691296022924,53.3900912448685 17.0553920767484,53.380195213511 17.0468579678559,53.3683369426613 17.0325277989031,53.3644639309539 17.0180045659715,53.2967628270739 16.9926640418376,53.2863539249682 16.9872160998117,53.2469410611709 16.9612614614385,53.1882110884165 16.9357962434572,53.158615811766 16.9251753342951,53.1437558398788 16.9208316662268,53.1471880142713 16.9142006024052,53.1380225074517 16.8974555042951,53.1295177539663 16.8610189642566,53.1327604006038 16.823481902673,53.1371541810432 16.7901437242966,53.1358036418982 16.7794762658421,53.1526103911524 16.7651159444561,53.1670519524728 16.7602795663432,53.1846195089798 16.7590843256964,53.1935880039937 16.76129287995,53.2036950623923 16.7556370018996,53.2381844323294 16.754214707265,53.2474508804875 16.7567061432602,53.2592756080982 16.74821459022,53.2651629915255 16.7500730986324,53.2907972143687 16.7493393703598,53.3080543225579 16.7468766614933,53.3162522784802 16.7411464199788,53.3320287901747 16.7427689590379,53.3390071658156 16.7388941275927,53.3474101380974 16.7423641283029,53.3697443313465 16.7352525259336,53.3961886814718 16.738457664686,53.4108890696058 16.7429642118719,53.4381114771362 16.7483901123903,53.4493847822058 16.7538052853579,53.4710396477033 16.7553409754229,53.4789246516732 16.7594199234924,53.5140938255255 16.7618497251788,53.518320872254 16.7594964572465,53.5501634493745 16.7582899312931,53.5593320691619 16.753765874908,53.5779444875584 16.7519098045522,53.5836709785499 16.7486861683579,53.589484635791 16.7545670217263,53.6093160480049 16.7616545267932,53.6415478396703 16.7706051496278,53.6570341916303 16.7780267638027,53.6741273481506 16.7826265023348,53.6706373535002 16.7940094479643,53.6752086813762 16.8058827871585,53.6866427877287 16.8164891888807,53.6907810011483 16.8150822347027,53.6999984260943 16.8240985692314,53.708843075719 16.8276607258778,53.7217395943175 16.8401013447786,53.7296343867967 16.8436002018834,53.7516462839885 16.8635340660338,53.754728287116 16.8702802043016))",Wilayat Rakhyut,ولاية رخيوت
"POLYGON ((55.6891378079147 18.9490818683714,55.0553759604434 19.9162032802052,55.0874155273192 19.961681388719,55.0573749325999 19.9984070021751,55.0102061953275 19.9845643688199,54.9999999983451 20.0000000436826,53.7610341920431 19.5941902700002,54.0462645146381 19.2764483805776,54.7725551691783 18.4590161358455,54.7824422325126 18.4629840636509,54.7872110223373 18.5003677105381,54.7853783843904 18.5219604618106,54.808825292255 18.5374924935908,54.81118371301 18.5567518641076,54.8560576436228 18.5969198042189,54.8784559444168 18.6124631062867,54.9086953521663 18.6596602408353,54.9546843242214 18.6997928398827,54.9518388834975 18.7214068071312,54.9759114607706 18.7766414513007,54.9921031628097 18.8002185110969,54.9975942516966 18.8160217276074,55.0001456251945 18.8443599826372,55.0277972884834 18.8563973757166,55.0661983983014 18.8784710557405,55.0781669397002 18.8987065213805,55.1166023246808 18.9219061973567,55.2287822075882 18.9256701840039,55.3579352899718 18.9313324723516,55.6891378079147 18.9490818683714))",Wilayat Muqshin,ولاية مقشن
"POLYGON ((56.5611249232296 24.5790028568444,56.5515917471391 24.5801493215928,56.5408350192318 24.563046489019,56.5105302293228 24.5508219456116,56.471676335606 24.5529461969283,56.4546593496852 24.5630348716339,56.4124642413297 24.5949702991384,56.4059805354049 24.6011696791035,56.3884509719013 24.6043321762625,56.3712525263257 24.5904284294458,56.3716645984331 24.5737554743686,56.3669107691476 24.539814788067,56.3135837026625 24.5498057807124,56.2753173397952 24.5464142738584,56.2376160493442 24.5408889023225,56.1940279816967 24.5362507248792,56.1969729975836 24.517662686419,56.2188323437681 24.4872011582328,56.2242442094765 24.4278873084447,56.2807538144619 24.4242911246786,56.342147885183 24.3758564884223,56.3260715090555 24.3381752190403,56.3526380889385 24.3372659420121,56.3607000680146 24.3290032358267,56.3667127733963 24.3104115843376,56.3866174562856 24.3117261954428,56.3899489261408 24.318397323314,56.40311480564 24.322518259343,56.4108570786259 24.3352569906318,56.4362030431712 24.3343753773861,56.4390051969048 24.3626835335924,56.4731402791766 24.3855327262649,56.4944876706013 24.3867425859019,56.529574454122 24.3967020543107,56.5339710064081 24.4048018244358,56.5344352864255 24.4179434524981,56.5427574436415 24.4315782992542,56.5594766838877 24.4388237198414,56.5662591564109 24.451680106998,56.5705506861093 24.4529307949604,56.6102078880428 24.4486008667109,56.6211558116319 24.454402267734,56.5837918629657 24.5114456638156,56.6032418590528 24.5227586929542,56.6000013592028 24.5308963306241,56.5927869659203 24.5359917616019,56.5611249232296 24.5790028568444))",Wilayat Liwa,ولاية لوى
"POLYGON ((56.1904192305869 26.2316974929453,56.1839382035111 26.2215228395501,56.184098447451 26.212212192413,56.1788309929929 26.2041684530167,56.1763892232796 26.1786717958141,56.1674184398008 26.1584415507903,56.1539194997211 26.1456320678166,56.141414206499 26.1453718825825,56.1308390767911 26.1273751774679,56.1249232073746 26.1126219832169,56.1127842182864 26.1018098080438,56.1019080768259 26.0863451471057,56.0988300313611 26.0756277707328,56.0902538925346 26.0677304148298,56.0861596801722 26.0554466830805,56.0894072279578 26.0509846177246,56.1070844506436 26.0556456681805,56.1165787453394 26.050593577435,56.1331824259423 26.0559401256501,56.1420086843952 26.0669813244879,56.1534079656728 26.0694232968556,56.1629263274727 26.0538402539497,56.1612788571849 26.0493612417794,56.1731005678016 26.0256012659566,56.1821800779531 26.0190886560574,56.1803761016021 25.9953675517307,56.1887316456723 25.9833063495997,56.1915264342557 25.9719811539477,56.1803468650122 25.9534713445222,56.1654631093071 25.9396075706244,56.1729009090257 25.9284718832061,56.1730978156654 25.9188567272974,56.1795793629032 25.9172050646558,56.1784278933725 25.89317130609,56.192628234753 25.8910078991936,56.1983194575243 25.8859230685461,56.2035814779468 25.8943376030323,56.1976818613242 25.9002216515776,56.1865286826783 25.9042710738121,56.2039079076113 25.9120499512568,56.2049656165275 25.9337376397275,56.2187358660179 25.935306449825,56.2216688500587 25.947674477187,56.1988108508504 25.9471154013325,56.1942910003635 25.9517605150518,56.192481341088 25.9632703048346,56.2005273739463 25.9826424682552,56.1995905899326 25.9963653951895,56.2081949619902 26.0041665919043,56.1835054493645 26.0387884390198,56.1780989220629 26.0493073597506,56.1880975403509 26.0549816947634,56.1781772328049 26.0721217043964,56.1739573703251 26.0867386066117,56.1841047380961 26.1182094777469,56.1961686112741 26.1341711141029,56.1869751838644 26.1462693583752,56.1928699651847 26.15914417088,56.1952471197256 26.176317285157,56.2024776643438 26.2051378571106,56.195238159047 26.2110917272221,56.202967093697 26.2206630534322,56.1904192305869 26.2316974929453))",Wilayat Bukha,ولاية بخاء
"MULTIPOLYGON (((56.4251519045391 25.9296128209767,56.4329749053474 25.9357364252369,56.4249545835743 25.9435008786837,56.4249503126604 25.9631586694512,56.4140267592646 25.9620650539769,56.4029076867093 25.9668825020856,56.4080229748585 25.9826373415982,56.4191610410089 25.9828783195759,56.4186450681845 25.9888017356404,56.4277887470465 25.9996654795807,56.4215867152315 26.0050842867664,56.4266601735747 26.0191079927335,56.4082134032272 26.0216788525752,56.4029642802066 26.0268553843742,56.39059355485 26.0174013141626,56.3873882526095 26.0338436853786,56.3905642192123 26.042229806767,56.405190251859 26.0456288104141,56.4170836723888 26.0414582538065,56.4367969365047 26.0434055669666,56.4356608482717 26.0591960310294,56.448359236664 26.071188900908,56.4583994862826 26.0738206515865,56.468564266451 26.0828811853844,56.4507166322464 26.0883155743481,56.4385413741776 26.0860248821056,56.43406267049 26.0895943458671,56.4173897730171 26.0806836188206,56.4092460577181 26.087849247806,56.4122417173721 26.0982476080278,56.3972884480597 26.0985109606807,56.390431848464 26.1044528506277,56.3788320838724 26.0869088661394,56.3700652348451 26.1081097131809,56.3790507129395 26.1272193052212,56.3612285685805 26.1251560315308,56.3470871186748 26.1090931053264,56.3469650549269 26.1001183534788,56.3336444885598 26.0957482551439,56.3369245553982 26.1061249238403,56.3355646520983 26.1179755501993,56.3390368735574 26.1250004454594,56.3331001428527 26.1419221203208,56.3354827452121 26.1494420016345,56.3266263128325 26.1539552313498,56.3331231171669 26.1651766269555,56.3432190703145 26.162061699007,56.3586476310986 26.1692860670825,56.3544547483802 26.1769110734089,56.3618361042072 26.1978223382832,56.3701087978693 26.1978429981051,56.3783956253191 26.2033327317756,56.3937260476903 26.1975133217107,56.3980910035615 26.1912021037345,56.3926780537314 26.1840439426269,56.3842132153505 26.1860124771263,56.3772781631607 26.1761926075965,56.3828504170097 26.168828364197,56.3785899071332 26.1580989949509,56.3826797705043 26.1528344186843,56.3926998171072 26.1798453999194,56.3987231918301 26.177443665027,56.4084476223931 26.1887922090059,56.4189389484799 26.1845611000088,56.4081398178973 26.1644330258003,56.414538130623 26.1637819819024,56.4150190933839 26.1529732485656,56.4197708182366 26.1397813199696,56.4300497539928 26.131596550483,56.4352021385357 26.1378019889663,56.4527298991973 26.1384475119248,56.4735828419935 26.1358976354121,56.4852123554395 26.1373708216571,56.4837609625645 26.146593734958,56.4719601741337 26.1426186391583,56.4735328061982 26.1517211242805,56.45840496996 26.1668230293788,56.4512044697047 26.1566641400058,56.4415917944393 26.1609976883242,56.4420827309439 26.1738110283252,56.4394888000682 26.1898530900289,56.4466430993809 26.1946153274753,56.4422091614298 26.2036429040504,56.4581387322949 26.2179079557933,56.470320004 26.2138219663311,56.4727435647938 26.2050914428585,56.4656695966908 26.1990199949405,56.4830020242649 26.1915872778404,56.483211575422 26.2010824339787,56.4748783127054 26.2117082069509,56.4733215229605 26.2248095804365,56.4790771040691 26.2319434188904,56.4745864971296 26.236893207012,56.453981548578 26.243917946394,56.4600991438803 26.2344760843217,56.453867827396 26.2274751326493,56.4445122451067 26.2238546444261,56.4315849579678 26.2334250456641,56.4252176563305 26.23098050363,56.4226885572561 26.2468043842496,56.4104409017269 26.2431991049736,56.3947933082831 26.2590234282958,56.4108914214043 26.2697876602336,56.4024798713988 26.2796913595699,56.3955353595279 26.2814500657098,56.4012611712226 26.2909264629745,56.4188571977428 26.2936873401022,56.4228707052487 26.2884237049536,56.4327377574862 26.2874190871953,56.4239634108273 26.3083688293317,56.4332983047723 26.3046811965201,56.4382013824168 26.3107888791512,56.4565300465151 26.3117583615344,56.4683274659793 26.318395272116,56.4811121497598 26.3161794680137,56.4981684781328 26.3190777022698,56.5044974560754 26.3129306291394,56.5145796636334 26.309863553501,56.5214072604313 26.317554610458,56.5060478687194 26.3206040755935,56.5085010824622 26.333203791516,56.5042344442298 26.3385976089609,56.5040218149261 26.353066198933,56.4953569704074 26.3503002929179,56.4915137791648 26.3355326088015,56.4990934348799 26.3286308059662,56.491475406813 26.3203693219051,56.4727346092572 26.3259353252123,56.4670793033246 26.321149156301,56.4508045119177 26.326891623345,56.4394289915995 26.3284082893652,56.4367590304251 26.3418326027959,56.429791390425 26.3520852806959,56.4144271974752 26.3379268323973,56.4098831107795 26.3389091651957,56.4176990751001 26.3629264020864,56.41173894059 26.3722336313525,56.403455204613 26.3563064192516,56.3962093692261 26.3555133728835,56.3885910372044 26.3697304121786,56.3781992438125 26.3651710375022,56.3685821226179 26.3657408598814,56.3694682010924 26.3541117932902,56.3598661857067 26.3345791169589,56.366984817945 26.3324001365937,56.3626517961174 26.3159954434191,56.3516616967545 26.3200385305537,56.3418928745476 26.3099056305242,56.3369301485514 26.31678344249,56.328415827023 26.3116350525931,56.3230351993716 26.3027115868979,56.3358662696697 26.2970242818303,56.341335336072 26.2874673295402,56.3489777195911 26.2869446522368,56.3549582985192 26.2782615920464,56.3690887207509 26.2741218517261,56.3631962955003 26.2681879527642,56.3765438617359 26.2594593096289,56.3676853542336 26.2480566027086,56.3617403612923 26.2523415779192,56.3459047755691 26.2533232360648,56.3484790686939 26.2660390784924,56.3409007661348 26.2679770041129,56.3351620644912 26.2775046489138,56.3195454207739 26.2856932354345,56.3144428633126 26.2663919326917,56.3140682964582 26.2575672337438,56.3189415556035 26.2489176527932,56.3089880786496 26.2419527078327,56.3033585214968 26.2293024014906,56.3018988250424 26.2183892625608,56.3053978319788 26.2040132257619,56.3105985560384 26.1987663642955,56.3266569658757 26.2021529034286,56.3331894560468 26.2060694257026,56.3403286295811 26.2194735492806,56.3518581718571 26.218365551402,56.3633509115019 26.2342038870199,56.3761796604761 26.2359254073705,56.3819453221677 26.2334690831137,56.3887823020256 26.2422276191362,56.394618655533 26.2384477624824,56.3912864803809 26.2297224409141,56.406592338089 26.2332436654795,56.4124559191372 26.2206341611111,56.4037918950306 26.2181743998995,56.4159535076379 26.2087730712364,56.3921689316953 26.2002052475664,56.3908341231529 26.2069715707042,56.3590534795691 26.2075281285975,56.3444244800166 26.1804656199435,56.3274024722191 26.1870224666788,56.3058794430452 26.1926569905195,56.2998152365768 26.1829400753468,56.2921656959852 26.1937210167341,56.2924852288977 26.2033485913241,56.2824533818639 26.2049096653104,56.2765132250097 26.2128953288673,56.2617129500895 26.2167683695637,56.2539501011844 26.2078264997494,56.2349170201915 26.2143901429884,56.2283551222778 26.2077107800315,56.2189372645692 26.2314030255491,56.218878478263 26.2521650553756,56.2076062254583 26.2529672649254,56.2057536117196 26.2451556974501,56.1959286143112 26.2402418830168,56.1904192305869 26.2316974929453,56.202967093697 26.2206630534322,56.195238159047 26.2110917272221,56.2024776643438 26.2051378571106,56.1952471197256 26.176317285157,56.1928699651847 26.15914417088,56.1869751838644 26.1462693583752,56.1961686112741 26.1341711141029,56.1841047380961 26.1182094777469,56.1739573703251 26.0867386066117,56.1781772328049 26.0721217043964,56.1880975403509 26.0549816947634,56.1780989220629 26.0493073597506,56.1835054493645 26.0387884390198,56.2081949619902 26.0041665919043,56.1995905899326 25.9963653951895,56.2005273739463 25.9826424682552,56.192481341088 25.9632703048346,56.1942910003635 25.9517605150518,56.1988108508504 25.9471154013325,56.2216688500587 25.947674477187,56.2187358660179 25.935306449825,56.2049656165275 25.9337376397275,56.2039079076113 25.9120499512568,56.1865286826783 25.9042710738121,56.1976818613242 25.9002216515776,56.2035814779468 25.8943376030323,56.1983194575243 25.8859230685461,56.2039551728054 25.8756452821828,56.2204107418475 25.8671836549533,56.2289421983578 25.8777155637139,56.2301632152982 25.8628697908512,56.2363265904557 25.8606865431743,56.2616285010419 25.8597061412811,56.2636878714708 25.8535643079505,56.2798420399877 25.8552601978985,56.2804926950215 25.8412040210082,56.2986293043029 25.8475115662234,56.310777736977 25.8642006006702,56.3160189954004 25.8839122131211,56.3261930340355 25.8916192868664,56.3349562960548 25.9030571080117,56.3359559583236 25.9139989377279,56.3491028255415 25.917920976859,56.3571379171061 25.9131041151726,56.3645616141125 25.9153620235197,56.3711245865737 25.9323467576518,56.3765818857828 25.9400710405254,56.3947859069078 25.9472857986561,56.4020221364435 25.9461760032619,56.4118504363211 25.9377984879004,56.4217143512012 25.9367509632418,56.4251519045391 25.9296128209767)),((56.3560817502548 26.375066563422,56.3447810671446 26.3552877394075,56.3420899873661 26.3359975414476,56.348300722989 26.3315207633557,56.3557321288314 26.3369384957712,56.3585267548874 26.3541331932706,56.3572148501561 26.3617486558776,56.3614497521197 26.3688652532709,56.3560817502548 26.375066563422)),((56.5266593059151 26.3875932960622,56.5222164133546 26.3678361985685,56.533496478317 26.3675438214359,56.5350975237311 26.377065818221,56.5266593059151 26.3875932960622)))",Wilayat Khasab,ولاية خصب
"MULTIPOLYGON (((58.7366961758017 20.9716858835556,58.7726505963806 21.0783795826631,58.8203522081033 21.1484771149746,58.9113066781793 21.1726683136766,58.9876202022621 21.2300498668939,59.0199964638301 21.2643067708461,59.0336917217238 21.2830373958973,58.9763343375928 21.2987081929137,58.9688792567802 21.3148045828243,58.9708013461071 21.3231995073333,58.9786721550959 21.3322057235353,58.9990780844017 21.3322636102079,59.0377677446359 21.3349484581808,59.0849490585331 21.3438158781291,59.2052519175106 21.415781910439,59.2403359439641 21.4426818720213,59.2445986161832 21.4535418106454,59.2577805667232 21.4743387452659,59.2571968518052 21.4769991642926,59.272307009337 21.505121193385,59.2751298305098 21.5456424560951,59.2576432383956 21.572961167066,59.2473636107754 21.5764666208211,59.2383411352088 21.5750075511621,59.2250956539978 21.5806406246003,59.1931691790532 21.6010088580843,59.1749684921411 21.6339453665669,59.1752751205448 21.6544082680953,59.2125107234575 21.66651304944,59.2494830933009 21.6612910939552,59.263633112307 21.6676656282726,59.2704572264111 21.6766813186801,59.2870791773548 21.7619519081237,59.2876678392423 21.7990484649778,59.2823257995707 21.8536224208283,59.2558435735687 21.907324952379,59.254398953735 21.9332015336058,59.2569188722626 21.9499119638339,59.2719545044043 21.9629552142052,59.2669152463076 21.970014212681,59.2570779326353 21.9698585896596,59.2310524004413 21.9527408475912,59.2175499186554 21.9476816164137,59.2098146714891 21.9521543351106,59.2117559482254 21.9692407970845,59.2100409540596 21.986664211126,59.228471805024 21.9980175688069,59.2484297430508 21.9967989545244,59.2616549564621 22.014719391487,59.277803641555 22.0254535814637,59.2847505185452 22.0267642274793,59.2851588405814 22.0382162913686,59.2916280114146 22.0428368958798,59.3042320411142 22.0434290087628,59.3165102584095 22.0571265182572,59.324208954164 22.0578949048719,59.3308747201718 22.0638809875231,59.3567964875126 22.0606486671379,59.3998872173722 22.0657807106554,59.4127104564645 22.0701978838535,59.4108535489606 22.1032816316995,59.4118880387445 22.1176576532123,59.4261958319379 22.1251826007808,59.4676571066379 22.1517449089695,59.4846353173464 22.1762019551284,59.4740102905363 22.2006633615444,59.4755842401944 22.2074151487596,59.4921926447481 22.2065160691032,59.5284380625384 22.2077387552054,59.5441351084601 22.2136679050294,59.5519151226396 22.2204718358326,59.5486036853776 22.2366888872238,59.5522234586209 22.2419328688639,59.5777099755223 22.2471363312277,59.6151298746662 22.2732768004873,59.6378774948486 22.2733074820527,59.6605145307538 22.2780438503401,59.7122808726534 22.3076848201277,59.7088911805478 22.3310394039781,59.6985990644119 22.3506996834679,59.6942466208153 22.3646565192907,59.6799520152513 22.399235125303,59.6540143480354 22.40734689121,59.6181154114187 22.4216904674893,59.5622919408316 22.4260255689457,59.5450109484815 22.4251524009108,59.5358171966832 22.416889168649,59.522260247519 22.3942857194129,59.5173877139838 22.3741910783058,59.5135826083804 22.3681812260475,59.5041278906553 22.3644909618743,59.4875470243662 22.3710483367528,59.4759486594778 22.3665677727163,59.4685299698081 22.3680940471434,59.454274869822 22.3602735525023,59.4463907405527 22.3711975231957,59.4292494145712 22.3652736923223,59.42192239865 22.3588808371624,59.4192415029776 22.3481635810561,59.4051327308771 22.3443628964766,59.3978379964327 22.3450805164122,59.3817720073295 22.3571270516784,59.3735038181256 22.3676066071158,59.363677211843 22.385906560427,59.3521537089643 22.3815539082376,59.3449064622558 22.3865278091828,59.328521746056 22.3882097102626,59.3180824112286 22.3651757600971,59.3182287640147 22.3557509258289,59.331803076603 22.3477988559574,59.343344014509 22.3346578633936,59.3433057583592 22.3265618482268,59.3561132838648 22.318257011333,59.3654952130732 22.3075770758188,59.3619937490122 22.2953287346222,59.3723040386607 22.2732994674986,59.3601192029617 22.2615139640533,59.3361026369146 22.2609335141734,59.3298661263579 22.2542333590579,59.3321725489509 22.2369168990017,59.3269375799301 22.2308584965844,59.3144777249982 22.2290339600684,59.3044401767764 22.2164279735702,59.3015387876658 22.201413034494,59.2894572809357 22.2004706007885,59.2808465370564 22.1787498499918,59.2704260923883 22.1446809004468,59.2580142259424 22.1350736069301,59.2451422807889 22.1509835288419,59.2389374010541 22.1541243755708,59.2310256614561 22.1496129056054,59.2158601768061 22.1720611443688,59.2106562390264 22.1760037594312,59.1969303456648 22.1755441300137,59.1856856200291 22.1696004975564,59.1669401856022 22.1698508772806,59.1600213253434 22.1862078935266,59.1375507972597 22.195578730064,59.1318951114234 22.2027054855092,59.1297383445964 22.2218177785633,59.1444649493334 22.2551908122804,59.1452985123342 22.2647310076705,59.1383302330333 22.2802186423179,59.1230013385636 22.2858527245142,59.0904368161967 22.2922986610043,59.0837304493275 22.297115514141,59.0887532777067 22.3229585335157,59.0798828581025 22.328090374862,59.0712199582506 22.3401651248328,59.0631964949916 22.3449178719158,59.0517012801913 22.3584025638822,59.0263228868264 22.3681118687284,59.0162964031917 22.3805023218107,59.0034754767876 22.3809426214505,59.0007021306189 22.3777937487495,59.0007620171919 22.3612699594903,59.0118048317269 22.3501207717276,59.0126037496748 22.2259469977024,59.0168293845203 22.2071179919954,59.0417927325163 22.1760867721844,59.0533764143827 22.1421999900346,59.0430958301371 22.126957993053,59.0365995639761 22.1214654755141,59.0340052142756 22.1053510244001,59.0130992180397 22.0757031128032,59.0063852256435 21.9605942956779,59.0080564118485 21.8946637595807,59.003217761385 21.8092019608218,58.9967498416596 21.6864656094361,58.9161844493334 21.658065424624,58.8954042203704 21.6187097107752,58.8859267519012 21.6062946274745,58.8688836672235 21.5939640265429,58.8480488999374 21.5935700156607,58.802488266457 21.6148680261066,58.7950775911053 21.6760432506166,58.8024397967133 21.7205115184638,58.7280327803024 21.7990127683807,58.7163255588312 21.7600806259773,58.7095299995633 21.7425158776126,58.7049853236941 21.7126196091186,58.7088867070958 21.6858177267404,58.7180354522144 21.668034601832,58.7438856506011 21.6444171127965,58.7561279649038 21.6287149562157,58.7596291065092 21.616457823968,58.7488949047067 21.5701763461444,58.7490444530929 21.5124175651795,58.7476758227008 21.4896644423517,58.7375137006501 21.4524385866533,58.6957080005763 21.3562265299308,58.6585153104252 21.204578716577,58.6497504597906 21.1833056833963,58.6452329337226 21.1623014932441,58.6395427210644 21.1585215313656,58.5868255477367 21.030369698721,58.6267497461294 21.0309071231811,58.6349361204547 20.9729287941786,58.7366961758017 20.9716858835556)),((59.3419779240712 21.4569056608148,59.3406392615121 21.4412027631222,59.3335177082995 21.435379622278,59.3126627505911 21.4352266158384,59.3054853765054 21.4453183818332,59.2988522942195 21.4606185922988,59.2893576224467 21.4528518816565,59.2895670993758 21.4395898689554,59.2847994904197 21.4276632647131,59.2891049285536 21.4233147156109,59.3064748045946 21.4263543815851,59.2982748941308 21.4140775158998,59.2994928296102 21.4097211776973,59.3436857427496 21.4329555220715,59.3514360095537 21.4449007154436,59.3419779240712 21.4569056608148)),((58.8642511792479 21.0768367784424,58.8555298407118 21.0811655141048,58.8315697311502 21.047196261012,58.8377470871983 21.0419754125787,58.8525507488148 21.0635125907971,58.8642511792479 21.0768367784424)),((59.1266189516903 21.319634815019,59.1134695894126 21.3191322234391,59.1048265563451 21.3244861476205,59.1042333005722 21.3138118499852,59.112348342781 21.3091017444302,59.1266189516903 21.319634815019)),((58.9450879610454 21.156961044257,58.9435489146352 21.166446597102,58.9359476114182 21.1632601635444,58.9310897325139 21.1479452798178,58.9214471207734 21.1393135656302,58.9450879610454 21.156961044257)),((59.0156552093212 21.2316408356765,59.029203241875 21.2454714187237,59.0123595036668 21.2391093327021,59.0156552093212 21.2316408356765)))",Wilayat Jaalan Bani Bu Hasan,ولاية جعلان بني بوحسن